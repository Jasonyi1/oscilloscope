
//
// Verific Verilog Description of module T35_Sensor_DDR3_LCD_Test
//

module T35_Sensor_DDR3_LCD_Test (clk_12M_i, Axi_Clk, tx_slowclk, tx_fastclk, 
            PllLocked, DdrCtrl_CFG_RST_N, DdrCtrl_CFG_SEQ_RST, DdrCtrl_CFG_SEQ_START, 
            DdrCtrl_AID_0, DdrCtrl_AADDR_0, DdrCtrl_ALEN_0, DdrCtrl_ASIZE_0, 
            DdrCtrl_ABURST_0, DdrCtrl_ALOCK_0, DdrCtrl_AVALID_0, DdrCtrl_AREADY_0, 
            DdrCtrl_ATYPE_0, DdrCtrl_WID_0, DdrCtrl_WDATA_0, DdrCtrl_WSTRB_0, 
            DdrCtrl_WLAST_0, DdrCtrl_WVALID_0, DdrCtrl_WREADY_0, DdrCtrl_RID_0, 
            DdrCtrl_RDATA_0, DdrCtrl_RLAST_0, DdrCtrl_RVALID_0, DdrCtrl_RREADY_0, 
            DdrCtrl_RRESP_0, DdrCtrl_BID_0, DdrCtrl_BVALID_0, DdrCtrl_BREADY_0, 
            LED, cmos_pclk, lcd_pwm, lvds_tx_clk_DATA, lvds_tx0_DATA, 
            lvds_tx1_DATA, lvds_tx2_DATA, lvds_tx3_DATA);
    input clk_12M_i /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input Axi_Clk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input tx_slowclk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input tx_fastclk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [1:0]PllLocked /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output DdrCtrl_CFG_RST_N /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_CFG_SEQ_RST /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_CFG_SEQ_START /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [7:0]DdrCtrl_AID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [31:0]DdrCtrl_AADDR_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [7:0]DdrCtrl_ALEN_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [2:0]DdrCtrl_ASIZE_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [1:0]DdrCtrl_ABURST_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [1:0]DdrCtrl_ALOCK_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_AVALID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input DdrCtrl_AREADY_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output DdrCtrl_ATYPE_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [7:0]DdrCtrl_WID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [127:0]DdrCtrl_WDATA_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [15:0]DdrCtrl_WSTRB_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_WLAST_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output DdrCtrl_WVALID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input DdrCtrl_WREADY_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]DdrCtrl_RID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [127:0]DdrCtrl_RDATA_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input DdrCtrl_RLAST_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input DdrCtrl_RVALID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output DdrCtrl_RREADY_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input [1:0]DdrCtrl_RRESP_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [7:0]DdrCtrl_BID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input DdrCtrl_BVALID_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output DdrCtrl_BREADY_0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [7:0]LED /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input cmos_pclk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output lcd_pwm /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx_clk_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx0_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx1_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx2_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [6:0]lvds_tx3_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]  /* verific async_reg="true" */ ;
    wire n6_2;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]  /* verific async_reg="true" */ ;
    wire \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]  /* verific async_reg="true" */ ;
    
    wire \ResetShiftReg[1] , n162, n163, \Axi0ResetReg[0] , \PowerOnResetCnt[0] , 
        \Axi0ResetReg[1] , \Axi0ResetReg[2] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0] , n176, n177, \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17] , \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19] , n198, n199, n200, 
        n201, \u_VsyHsyGenerator/pCnt_value[0] , \u_VsyHsyGenerator/frameCnt_value[0] , 
        \u_VsyHsyGenerator/vsynDl[0] , \u_VsyHsyGenerator/pCntInc , \u_VsyHsyGenerator/hsynDl[0] , 
        \u_VsyHsyGenerator/hsynCnt_value[0] , n216, n217, n218, n219, 
        n220, n221, n222, n223, n224, n225, n226, n227, n228, 
        n229, n230, n231, n232, n233, n234, n235, n236, n237, 
        n238, n239, n240, n241, n242, n243, n244, n245, n246, 
        n247, n248, n249, n250, n251, n252, n253, n254, n255, 
        n256, n257, n258, n259, n260, n261, n262, n263, n264, 
        n265, n266, n267, n268, n269, n270, n271, n272, n273, 
        n274, n275, n276, n277, n278, n279, n280, n281, n282, 
        n283, n284, n285, n286, n287, n288, n289, n290, n291, 
        n292, n293, n294, n295, n296, n297, n298, n299, n300, 
        n301, n303, n305, n307, n309, n311, n312, n313, n314, 
        n315, n316, n317, n318, n319, n320, n321, n322, n323, 
        n324, n325, n326, n327, n328, n329, n330, n331, n332, 
        n333, n334, n335, n336, n337, n338, n339, n340, n341, 
        n342, n343, n344, n345, \u_VsyHsyGenerator/pCnt_value[1] , 
        \u_VsyHsyGenerator/pCnt_value[2] , \u_VsyHsyGenerator/pCnt_value[3] , 
        \u_VsyHsyGenerator/pCnt_value[4] , \u_VsyHsyGenerator/pCnt_value[5] , 
        \u_VsyHsyGenerator/pCnt_value[6] , \u_VsyHsyGenerator/pCnt_value[7] , 
        \u_VsyHsyGenerator/pCnt_value[8] , \u_VsyHsyGenerator/pCnt_value[9] , 
        \u_VsyHsyGenerator/pCnt_value[10] , \u_VsyHsyGenerator/frameCnt_value[1] , 
        \u_VsyHsyGenerator/frameCnt_value[2] , \u_VsyHsyGenerator/frameCnt_value[3] , 
        \u_VsyHsyGenerator/frameCnt_value[4] , \u_VsyHsyGenerator/frameCnt_value[5] , 
        \u_VsyHsyGenerator/frameCnt_value[6] , \u_VsyHsyGenerator/frameCnt_value[7] , 
        \u_VsyHsyGenerator/frameCnt_value[8] , \u_VsyHsyGenerator/frameCnt_value[9] , 
        \u_VsyHsyGenerator/vsynDl[1] , \u_VsyHsyGenerator/vsynDl[2] , XYCrop_frame_vsync, 
        \u_VsyHsyGenerator/hsynDl[1] , \u_VsyHsyGenerator/hsynDl[2] , XYCrop_frame_href, 
        \u_VsyHsyGenerator/hsynCnt_value[1] , \u_VsyHsyGenerator/hsynCnt_value[2] , 
        \u_VsyHsyGenerator/hsynCnt_value[3] , \u_VsyHsyGenerator/hsynCnt_value[4] , 
        \u_VsyHsyGenerator/hsynCnt_value[5] , \u_VsyHsyGenerator/hsynCnt_value[6] , 
        \u_VsyHsyGenerator/hsynCnt_value[7] , \u_VsyHsyGenerator/hsynCnt_value[8] , 
        \u_VsyHsyGenerator/hsynCnt_value[9] , n380, n381, n382, \u_axi4_ctrl/wframe_vsync_dly[0] , 
        \u_axi4_ctrl/wframe_index[1] , \u_axi4_ctrl/rframe_vsync_dly[0] , 
        \u_axi4_ctrl/wfifo_cnt[0] , \u_axi4_ctrl/wfifo_rst , \u_axi4_ctrl/wframe_index[0] , 
        n397, n398, n399, n400, n401, n402, \u_axi4_ctrl/rframe_index[0] , 
        \u_axi4_ctrl/state[0] , n405, n406, \u_axi4_ctrl/wframe_vsync_dly[1] , 
        n409, n410, n411, n412, n413, n414, n415, n416, n418, 
        n419, n420, n421, n422, n423, \u_axi4_ctrl/wframe_vsync_dly[3] , 
        n425, n426, n427, n460, n461, n470, n471, n480, n481, 
        n482, n483, n484, n485, n486, n487, n488, n489, n490, 
        n491, n516, n517, \u_axi4_ctrl/wfifo_cnt[4] , \u_axi4_ctrl/wfifo_cnt[3] , 
        n539, n540, n541, n542, n543, n544, \u_axi4_ctrl/wdata_cnt_dly[0] , 
        \u_axi4_ctrl/rdata_cnt_dly[1] , \u_axi4_ctrl/rdata_cnt_dly[0] , 
        \u_axi4_ctrl/wfifo_cnt[2] , \u_axi4_ctrl/wfifo_cnt[1] , \u_axi4_ctrl/rframe_vsync_dly[3] , 
        n551, n552, n553, n554, n555, \u_axi4_ctrl/rfifo_wenb , 
        n559, n560, \u_axi4_ctrl/rfifo_wdata[0] , n563, n564, n565, 
        n566, \lcd_data[0] , \lcd_data[1] , n569, n570, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/wfifo_empty , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12] , 
        n593, n594, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , 
        n597, n598, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
        n601, n602, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
        n613, \lcd_data[4] , \lcd_data[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[9] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12] , 
        n713, n714, n715, n716, n717, n718, n719, n720, n721, 
        n722, n723, n724, n725, n726, n727, n728, \lcd_data[6] , 
        \lcd_data[7] , \lcd_data[10] , \lcd_data[11] , \lcd_data[12] , 
        \lcd_data[13] , \lcd_data[14] , \lcd_data[15] , \lcd_data[8] , 
        \lcd_data[9] , n747, n748, \lcd_data[2] , \lcd_data[3] , n754, 
        n755, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] , \u_axi4_ctrl/rfifo_empty , 
        n758, n759, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] , n761, 
        n762, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] , 
        n766, n767, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] , 
        n776, n777, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[11] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] , 
        n869, n870, \u_axi4_ctrl/rframe_index[1] , \u_axi4_ctrl/state[1] , 
        \u_axi4_ctrl/state[2] , \u_axi4_ctrl/awaddr[10] , \u_axi4_ctrl/awaddr[11] , 
        \u_axi4_ctrl/awaddr[12] , \u_axi4_ctrl/awaddr[13] , \u_axi4_ctrl/awaddr[14] , 
        \u_axi4_ctrl/awaddr[15] , \u_axi4_ctrl/awaddr[16] , \u_axi4_ctrl/awaddr[17] , 
        \u_axi4_ctrl/awaddr[18] , \u_axi4_ctrl/awaddr[19] , \u_axi4_ctrl/awaddr[20] , 
        \u_axi4_ctrl/awaddr[21] , \u_axi4_ctrl/awaddr[22] , \u_axi4_ctrl/awaddr[23] , 
        n888, n889, n890, n891, n892, n893, n894, n895, n896, 
        n897, n898, n899, n900, n901, n902, n903, n904, n905, 
        n906, n907, n908, n909, n910, n911, n912, n913, n914, 
        n915, n916, n917, n918, n919, n920, n921, n922, n923, 
        n924, n925, n926, n927, n928, n929, n930, n931, \u_axi4_ctrl/araddr[10] , 
        \u_axi4_ctrl/araddr[11] , \u_axi4_ctrl/araddr[12] , \u_axi4_ctrl/araddr[13] , 
        \u_axi4_ctrl/araddr[14] , \u_axi4_ctrl/araddr[15] , \u_axi4_ctrl/araddr[16] , 
        \u_axi4_ctrl/araddr[17] , \u_axi4_ctrl/araddr[18] , \u_axi4_ctrl/araddr[19] , 
        \u_axi4_ctrl/araddr[20] , \u_axi4_ctrl/araddr[21] , \u_axi4_ctrl/araddr[22] , 
        \u_axi4_ctrl/araddr[23] , n946, n947, n948, n949, n950, 
        n951, n952, n953, n954, n955, n956, n957, n958, n959, 
        n960, n961, n962, n963, n964, n965, n966, n967, n968, 
        n969, n970, n971, n972, n989, n990, \u_axi4_ctrl/wdata_cnt_dly[1] , 
        \u_axi4_ctrl/wdata_cnt_dly[2] , \u_axi4_ctrl/wdata_cnt_dly[3] , 
        \u_axi4_ctrl/wdata_cnt_dly[4] , \u_axi4_ctrl/wdata_cnt_dly[5] , 
        \u_axi4_ctrl/wdata_cnt_dly[6] , \u_axi4_ctrl/wdata_cnt_dly[7] , 
        \u_axi4_ctrl/wdata_cnt_dly[8] , \u_axi4_ctrl/rdata_cnt_dly[2] , 
        \u_axi4_ctrl/rdata_cnt_dly[3] , \u_axi4_ctrl/rdata_cnt_dly[4] , 
        \u_axi4_ctrl/rdata_cnt_dly[5] , \u_axi4_ctrl/rdata_cnt_dly[6] , 
        \u_axi4_ctrl/rdata_cnt_dly[7] , \u_axi4_ctrl/rdata_cnt_dly[8] , 
        n1006, n1007, n1008, n1009, \u_axi4_ctrl/rfifo_wdata[1] , 
        \u_axi4_ctrl/rfifo_wdata[2] , \u_axi4_ctrl/rfifo_wdata[3] , \u_axi4_ctrl/rfifo_wdata[4] , 
        \u_axi4_ctrl/rfifo_wdata[5] , \u_axi4_ctrl/rfifo_wdata[6] , \u_axi4_ctrl/rfifo_wdata[7] , 
        \u_axi4_ctrl/rfifo_wdata[8] , \u_axi4_ctrl/rfifo_wdata[9] , \u_axi4_ctrl/rfifo_wdata[10] , 
        \u_axi4_ctrl/rfifo_wdata[11] , \u_axi4_ctrl/rfifo_wdata[12] , \u_axi4_ctrl/rfifo_wdata[13] , 
        \u_axi4_ctrl/rfifo_wdata[14] , \u_axi4_ctrl/rfifo_wdata[15] , \u_axi4_ctrl/rfifo_wdata[16] , 
        \u_axi4_ctrl/rfifo_wdata[17] , \u_axi4_ctrl/rfifo_wdata[18] , \u_axi4_ctrl/rfifo_wdata[19] , 
        \u_axi4_ctrl/rfifo_wdata[20] , \u_axi4_ctrl/rfifo_wdata[21] , \u_axi4_ctrl/rfifo_wdata[22] , 
        \u_axi4_ctrl/rfifo_wdata[23] , \u_axi4_ctrl/rfifo_wdata[24] , \u_axi4_ctrl/rfifo_wdata[25] , 
        \u_axi4_ctrl/rfifo_wdata[26] , \u_axi4_ctrl/rfifo_wdata[27] , \u_axi4_ctrl/rfifo_wdata[28] , 
        \u_axi4_ctrl/rfifo_wdata[29] , \u_axi4_ctrl/rfifo_wdata[30] , \u_axi4_ctrl/rfifo_wdata[31] , 
        \u_axi4_ctrl/rfifo_wdata[32] , \u_axi4_ctrl/rfifo_wdata[33] , \u_axi4_ctrl/rfifo_wdata[34] , 
        \u_axi4_ctrl/rfifo_wdata[35] , \u_axi4_ctrl/rfifo_wdata[36] , \u_axi4_ctrl/rfifo_wdata[37] , 
        \u_axi4_ctrl/rfifo_wdata[38] , \u_axi4_ctrl/rfifo_wdata[39] , \u_axi4_ctrl/rfifo_wdata[40] , 
        \u_axi4_ctrl/rfifo_wdata[41] , \u_axi4_ctrl/rfifo_wdata[42] , \u_axi4_ctrl/rfifo_wdata[43] , 
        \u_axi4_ctrl/rfifo_wdata[44] , \u_axi4_ctrl/rfifo_wdata[45] , \u_axi4_ctrl/rfifo_wdata[46] , 
        \u_axi4_ctrl/rfifo_wdata[47] , \u_axi4_ctrl/rfifo_wdata[48] , \u_axi4_ctrl/rfifo_wdata[49] , 
        \u_axi4_ctrl/rfifo_wdata[50] , \u_axi4_ctrl/rfifo_wdata[51] , \u_axi4_ctrl/rfifo_wdata[52] , 
        \u_axi4_ctrl/rfifo_wdata[53] , \u_axi4_ctrl/rfifo_wdata[54] , \u_axi4_ctrl/rfifo_wdata[55] , 
        \u_axi4_ctrl/rfifo_wdata[56] , \u_axi4_ctrl/rfifo_wdata[57] , \u_axi4_ctrl/rfifo_wdata[58] , 
        \u_axi4_ctrl/rfifo_wdata[59] , \u_axi4_ctrl/rfifo_wdata[60] , \u_axi4_ctrl/rfifo_wdata[61] , 
        \u_axi4_ctrl/rfifo_wdata[62] , \u_axi4_ctrl/rfifo_wdata[63] , \u_axi4_ctrl/rfifo_wdata[64] , 
        \u_axi4_ctrl/rfifo_wdata[65] , \u_axi4_ctrl/rfifo_wdata[66] , \u_axi4_ctrl/rfifo_wdata[67] , 
        \u_axi4_ctrl/rfifo_wdata[68] , \u_axi4_ctrl/rfifo_wdata[69] , \u_axi4_ctrl/rfifo_wdata[70] , 
        \u_axi4_ctrl/rfifo_wdata[71] , \u_axi4_ctrl/rfifo_wdata[72] , \u_axi4_ctrl/rfifo_wdata[73] , 
        \u_axi4_ctrl/rfifo_wdata[74] , \u_axi4_ctrl/rfifo_wdata[75] , \u_axi4_ctrl/rfifo_wdata[76] , 
        \u_axi4_ctrl/rfifo_wdata[77] , \u_axi4_ctrl/rfifo_wdata[78] , \u_axi4_ctrl/rfifo_wdata[79] , 
        \u_axi4_ctrl/rfifo_wdata[80] , \u_axi4_ctrl/rfifo_wdata[81] , \u_axi4_ctrl/rfifo_wdata[82] , 
        \u_axi4_ctrl/rfifo_wdata[83] , \u_axi4_ctrl/rfifo_wdata[84] , \u_axi4_ctrl/rfifo_wdata[85] , 
        \u_axi4_ctrl/rfifo_wdata[86] , \u_axi4_ctrl/rfifo_wdata[87] , \u_axi4_ctrl/rfifo_wdata[88] , 
        \u_axi4_ctrl/rfifo_wdata[89] , \u_axi4_ctrl/rfifo_wdata[90] , \u_axi4_ctrl/rfifo_wdata[91] , 
        \u_axi4_ctrl/rfifo_wdata[92] , \u_axi4_ctrl/rfifo_wdata[93] , \u_axi4_ctrl/rfifo_wdata[94] , 
        \u_axi4_ctrl/rfifo_wdata[95] , \u_axi4_ctrl/rfifo_wdata[96] , \u_axi4_ctrl/rfifo_wdata[97] , 
        \u_axi4_ctrl/rfifo_wdata[98] , \u_axi4_ctrl/rfifo_wdata[99] , \u_axi4_ctrl/rfifo_wdata[100] , 
        \u_axi4_ctrl/rfifo_wdata[101] , \u_axi4_ctrl/rfifo_wdata[102] , 
        \u_axi4_ctrl/rfifo_wdata[103] , \u_axi4_ctrl/rfifo_wdata[104] , 
        \u_axi4_ctrl/rfifo_wdata[105] , \u_axi4_ctrl/rfifo_wdata[106] , 
        \u_axi4_ctrl/rfifo_wdata[107] , \u_axi4_ctrl/rfifo_wdata[108] , 
        \u_axi4_ctrl/rfifo_wdata[109] , \u_axi4_ctrl/rfifo_wdata[110] , 
        \u_axi4_ctrl/rfifo_wdata[111] , \u_axi4_ctrl/rfifo_wdata[112] , 
        \u_axi4_ctrl/rfifo_wdata[113] , \u_axi4_ctrl/rfifo_wdata[114] , 
        \u_axi4_ctrl/rfifo_wdata[115] , \u_axi4_ctrl/rfifo_wdata[116] , 
        \u_axi4_ctrl/rfifo_wdata[117] , \u_axi4_ctrl/rfifo_wdata[118] , 
        \u_axi4_ctrl/rfifo_wdata[119] , \u_axi4_ctrl/rfifo_wdata[120] , 
        \u_axi4_ctrl/rfifo_wdata[121] , \u_axi4_ctrl/rfifo_wdata[122] , 
        \u_axi4_ctrl/rfifo_wdata[123] , \u_axi4_ctrl/rfifo_wdata[124] , 
        \u_axi4_ctrl/rfifo_wdata[125] , \u_axi4_ctrl/rfifo_wdata[126] , 
        \u_axi4_ctrl/rfifo_wdata[127] , n1137, n1138, \u_lcd_driver/vcnt[0] , 
        n1140, n1141, n1142, n1143, \u_lcd_driver/hcnt[0] , \u_lcd_driver/vcnt[1] , 
        \u_lcd_driver/vcnt[2] , \u_lcd_driver/vcnt[3] , \u_lcd_driver/vcnt[4] , 
        \u_lcd_driver/vcnt[5] , \u_lcd_driver/vcnt[6] , \u_lcd_driver/vcnt[7] , 
        \u_lcd_driver/vcnt[8] , \u_lcd_driver/vcnt[9] , \u_lcd_driver/vcnt[10] , 
        \u_lcd_driver/vcnt[11] , n1156, n1157, n1158, n1159, n1160, 
        n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, 
        n1169, n1170, n1171, n1172, n1173, n1174, \u_lcd_driver/hcnt[1] , 
        \u_lcd_driver/hcnt[2] , \u_lcd_driver/hcnt[3] , \u_lcd_driver/hcnt[4] , 
        \u_lcd_driver/hcnt[5] , \u_lcd_driver/hcnt[6] , \u_lcd_driver/hcnt[7] , 
        \u_lcd_driver/hcnt[8] , \u_lcd_driver/hcnt[9] , \u_lcd_driver/hcnt[10] , 
        \u_lcd_driver/hcnt[11] , \PowerOnResetCnt[1] , \PowerOnResetCnt[2] , 
        \PowerOnResetCnt[3] , \PowerOnResetCnt[4] , \PowerOnResetCnt[5] , 
        \PowerOnResetCnt[6] , \PowerOnResetCnt[7] , \ResetShiftReg[0] , 
        \reduce_nand_6/n7 , DdrInitDone, \U0_DDR_Reset/u_ddr_reset_sequencer/n15 , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/equal_21/n3 , \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] , 
        \U0_DDR_Reset/u_ddr_reset_sequencer/n92 , \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0] , 
        n1405, \U0_DDR_Reset/u_ddr_reset_sequencer/n91 , n1429, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int , 
        \XYCrop_frame_Gray[15] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int , 
        \u_VsyHsyGenerator/pCnt_valueNext[0] , \u_VsyHsyGenerator/frameCnt_valueNext[0] , 
        \u_VsyHsyGenerator/n402 , ceg_net2, \u_VsyHsyGenerator/when_MyTopLevel_l56 , 
        ceg_net5, \u_VsyHsyGenerator/n519 , \u_VsyHsyGenerator/hsynCnt_valueNext[0] , 
        n1553, n1556, n1559, n1562, n1565, n1568, n1571, n1574, 
        \u_VsyHsyGenerator/pCnt_valueNext[1] , \u_VsyHsyGenerator/pCnt_valueNext[2] , 
        \u_VsyHsyGenerator/pCnt_valueNext[3] , \u_VsyHsyGenerator/pCnt_valueNext[4] , 
        \u_VsyHsyGenerator/pCnt_valueNext[5] , \u_VsyHsyGenerator/pCnt_valueNext[6] , 
        \u_VsyHsyGenerator/pCnt_valueNext[7] , \u_VsyHsyGenerator/pCnt_valueNext[8] , 
        \u_VsyHsyGenerator/pCnt_valueNext[9] , \u_VsyHsyGenerator/pCnt_valueNext[10] , 
        \u_VsyHsyGenerator/frameCnt_valueNext[1] , \u_VsyHsyGenerator/frameCnt_valueNext[2] , 
        \u_VsyHsyGenerator/frameCnt_valueNext[3] , \u_VsyHsyGenerator/frameCnt_valueNext[4] , 
        \u_VsyHsyGenerator/frameCnt_valueNext[5] , \u_VsyHsyGenerator/frameCnt_valueNext[6] , 
        \u_VsyHsyGenerator/frameCnt_valueNext[7] , \u_VsyHsyGenerator/frameCnt_valueNext[8] , 
        \u_VsyHsyGenerator/frameCnt_valueNext[9] , \u_VsyHsyGenerator/n681 , 
        \u_VsyHsyGenerator/n416 , \u_VsyHsyGenerator/n415 , \u_VsyHsyGenerator/n414 , 
        \u_VsyHsyGenerator/hsynCnt_valueNext[1] , \u_VsyHsyGenerator/hsynCnt_valueNext[2] , 
        \u_VsyHsyGenerator/hsynCnt_valueNext[3] , \u_VsyHsyGenerator/hsynCnt_valueNext[4] , 
        \u_VsyHsyGenerator/hsynCnt_valueNext[5] , \u_VsyHsyGenerator/hsynCnt_valueNext[6] , 
        \u_VsyHsyGenerator/hsynCnt_valueNext[7] , \u_VsyHsyGenerator/hsynCnt_valueNext[8] , 
        \u_VsyHsyGenerator/hsynCnt_valueNext[9] , \u_axi4_ctrl/n323 , \u_axi4_ctrl/equal_37/n3 , 
        \u_lcd_driver/n108 , \u_axi4_ctrl/n96 , \u_axi4_ctrl/n1476 , \u_axi4_ctrl/equal_28/n9 , 
        \u_axi4_ctrl/n324 , \XYCrop_frame_Gray[14] , \u_axi4_ctrl/n343 , 
        \u_axi4_ctrl/equal_46/n3 , \u_axi4_ctrl/n396 , \u_axi4_ctrl/n412 , 
        \u_axi4_ctrl/n1483 , \u_axi4_ctrl/wframe_vsync_dly[2] , \XYCrop_frame_Gray[9] , 
        \XYCrop_frame_Gray[5] , \u_axi4_ctrl/n92 , \u_axi4_ctrl/n93 , 
        \u_axi4_ctrl/n370 , \u_axi4_ctrl/n1551 , \u_axi4_ctrl/n386 , \u_axi4_ctrl/n94 , 
        \u_axi4_ctrl/n95 , \u_axi4_ctrl/rframe_vsync_dly[2] , \u_axi4_ctrl/rframe_vsync_dly[1] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int , 
        ceg_net12, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[0] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] , 
        n1776, \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[1] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[9] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[10] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[11] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[9] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[8] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[9] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[10] , 
        \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[11] , 
        ceg_net19, \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[0] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[8] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[9] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[10] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[1] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[8] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[9] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[10] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[11] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] , 
        \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] , 
        \u_axi4_ctrl/n342 , \u_axi4_ctrl/n1616 , \u_axi4_ctrl/n1623 , 
        \u_axi4_ctrl/n394 , \u_axi4_ctrl/n376 , \u_axi4_ctrl/n388 , \u_axi4_ctrl/n1485 , 
        \u_axi4_ctrl/n704 , ceg_net124, \u_axi4_ctrl/n703 , \u_axi4_ctrl/n702 , 
        \u_axi4_ctrl/n701 , \u_axi4_ctrl/n700 , \u_axi4_ctrl/n699 , \u_axi4_ctrl/n698 , 
        \u_axi4_ctrl/n697 , \u_axi4_ctrl/n696 , \u_axi4_ctrl/n695 , \u_axi4_ctrl/n694 , 
        \u_axi4_ctrl/n693 , \u_axi4_ctrl/n692 , \u_axi4_ctrl/n691 , \u_axi4_ctrl/n690 , 
        \u_axi4_ctrl/n689 , \u_axi4_ctrl/n1506 , \u_axi4_ctrl/n1511 , 
        \u_axi4_ctrl/n1516 , \u_axi4_ctrl/n1521 , \u_axi4_ctrl/n1526 , 
        \u_axi4_ctrl/n1531 , \u_axi4_ctrl/n1536 , \u_axi4_ctrl/n1541 , 
        \u_axi4_ctrl/n1556 , \u_axi4_ctrl/n1561 , \u_axi4_ctrl/n1566 , 
        \u_axi4_ctrl/n1571 , \u_axi4_ctrl/n1576 , \u_axi4_ctrl/n1581 , 
        \u_axi4_ctrl/n1586 , \u_lcd_driver/n81 , \u_lcd_driver/equal_15/n23 , 
        \u_lcd_driver/n34 , \u_lcd_driver/n80 , \u_lcd_driver/n79 , \u_lcd_driver/n78 , 
        \u_lcd_driver/n77 , \u_lcd_driver/n76 , \u_lcd_driver/n75 , \u_lcd_driver/n74 , 
        \u_lcd_driver/n73 , \u_lcd_driver/n72 , \u_lcd_driver/n71 , \u_lcd_driver/n70 , 
        \tx_slowclk~O , \u_lcd_driver/n33 , \u_lcd_driver/n32 , \u_lcd_driver/n31 , 
        \u_lcd_driver/n30 , \u_lcd_driver/n29 , \u_lcd_driver/n28 , \u_lcd_driver/n27 , 
        \u_lcd_driver/n26 , \u_lcd_driver/n25 , \u_lcd_driver/n24 , \u_lcd_driver/n23 , 
        \clk_12M_i~O , \Axi_Clk~O , n2556, n2555, n2554, n2553, 
        n2552, n2429, n2430, n2431, n2432, n2433, n2434, n2435, 
        n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, 
        n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, 
        n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, 
        n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, 
        n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, 
        n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, 
        n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, 
        n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, 
        n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, 
        n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, 
        n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, 
        n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, 
        n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, 
        n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, 
        n2548, n2549, n2550, n2551;
    
    assign DdrCtrl_AID_0[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AID_0[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[31] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[30] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[29] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[28] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[27] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[26] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[9] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[8] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_AADDR_0[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[5] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[4] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[3] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[2] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[1] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALEN_0[0] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ASIZE_0[2] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ASIZE_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ASIZE_0[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ABURST_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALOCK_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_ALOCK_0[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WID_0[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[15] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[14] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[13] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[12] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[11] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[10] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[9] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[8] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[7] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[6] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[5] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[4] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[3] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[2] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[1] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign DdrCtrl_WSTRB_0[0] = DdrCtrl_ABURST_0[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign LED[7] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign LED[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign LED[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign LED[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign LED[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign LED[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign LED[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign LED[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lcd_pwm = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[6] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[5] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[0] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx0_DATA[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx1_DATA[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx2_DATA[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx3_DATA[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign lvds_tx_clk_DATA[1] = 1'b1 /* verific EFX_ATTRIBUTE_CELL_NAME=VCC */ ;
    assign DdrCtrl_WID_0[0] = 1'b0 /* verific EFX_ATTRIBUTE_CELL_NAME=GND */ ;
    EFX_LUT4 LUT__3686 (.I0(\u_axi4_ctrl/state[2] ), .I1(\u_axi4_ctrl/state[1] ), 
            .O(DdrCtrl_BREADY_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3686.LUTMASK = 16'h4444;
    EFX_FF \ResetShiftReg[1]~FF  (.D(\ResetShiftReg[0] ), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\ResetShiftReg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(106)
    defparam \ResetShiftReg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \ResetShiftReg[1]~FF .CE_POLARITY = 1'b1;
    defparam \ResetShiftReg[1]~FF .SR_POLARITY = 1'b1;
    defparam \ResetShiftReg[1]~FF .D_POLARITY = 1'b1;
    defparam \ResetShiftReg[1]~FF .SR_SYNC = 1'b1;
    defparam \ResetShiftReg[1]~FF .SR_VALUE = 1'b0;
    defparam \ResetShiftReg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \ResetShiftReg[0]~FF  (.D(\reduce_nand_6/n7 ), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\ResetShiftReg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(106)
    defparam \ResetShiftReg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \ResetShiftReg[0]~FF .CE_POLARITY = 1'b1;
    defparam \ResetShiftReg[0]~FF .SR_POLARITY = 1'b1;
    defparam \ResetShiftReg[0]~FF .D_POLARITY = 1'b1;
    defparam \ResetShiftReg[0]~FF .SR_SYNC = 1'b1;
    defparam \ResetShiftReg[0]~FF .SR_VALUE = 1'b0;
    defparam \ResetShiftReg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \Axi0ResetReg[0]~FF  (.D(DdrInitDone), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\Axi0ResetReg[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(139)
    defparam \Axi0ResetReg[0]~FF .CLK_POLARITY = 1'b1;
    defparam \Axi0ResetReg[0]~FF .CE_POLARITY = 1'b1;
    defparam \Axi0ResetReg[0]~FF .SR_POLARITY = 1'b1;
    defparam \Axi0ResetReg[0]~FF .D_POLARITY = 1'b1;
    defparam \Axi0ResetReg[0]~FF .SR_SYNC = 1'b1;
    defparam \Axi0ResetReg[0]~FF .SR_VALUE = 1'b0;
    defparam \Axi0ResetReg[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_CFG_RST_N~FF  (.D(\ResetShiftReg[1] ), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(DdrCtrl_CFG_RST_N)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(106)
    defparam \DdrCtrl_CFG_RST_N~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_RST_N~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_RST_N~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_RST_N~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_RST_N~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_CFG_RST_N~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_CFG_RST_N~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[0]~FF  (.D(n1173), .CE(n6_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(99)
    defparam \PowerOnResetCnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[0]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \Axi0ResetReg[1]~FF  (.D(\Axi0ResetReg[0] ), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\Axi0ResetReg[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(139)
    defparam \Axi0ResetReg[1]~FF .CLK_POLARITY = 1'b1;
    defparam \Axi0ResetReg[1]~FF .CE_POLARITY = 1'b1;
    defparam \Axi0ResetReg[1]~FF .SR_POLARITY = 1'b1;
    defparam \Axi0ResetReg[1]~FF .D_POLARITY = 1'b1;
    defparam \Axi0ResetReg[1]~FF .SR_SYNC = 1'b1;
    defparam \Axi0ResetReg[1]~FF .SR_VALUE = 1'b0;
    defparam \Axi0ResetReg[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \Axi0ResetReg[2]~FF  (.D(\Axi0ResetReg[1] ), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\Axi0ResetReg[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(139)
    defparam \Axi0ResetReg[2]~FF .CLK_POLARITY = 1'b1;
    defparam \Axi0ResetReg[2]~FF .CE_POLARITY = 1'b1;
    defparam \Axi0ResetReg[2]~FF .SR_POLARITY = 1'b1;
    defparam \Axi0ResetReg[2]~FF .D_POLARITY = 1'b1;
    defparam \Axi0ResetReg[2]~FF .SR_SYNC = 1'b1;
    defparam \Axi0ResetReg[2]~FF .SR_VALUE = 1'b0;
    defparam \Axi0ResetReg[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrInitDone~FF  (.D(1'b1), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(DdrInitDone)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \DdrInitDone~FF .CLK_POLARITY = 1'b1;
    defparam \DdrInitDone~FF .CE_POLARITY = 1'b0;
    defparam \DdrInitDone~FF .SR_POLARITY = 1'b0;
    defparam \DdrInitDone~FF .D_POLARITY = 1'b1;
    defparam \DdrInitDone~FF .SR_SYNC = 1'b0;
    defparam \DdrInitDone~FF .SR_VALUE = 1'b0;
    defparam \DdrInitDone~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_CFG_SEQ_START~FF  (.D(1'b1), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/equal_21/n3 ), 
           .CLK(\Axi_Clk~O ), .SR(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] ), 
           .Q(DdrCtrl_CFG_SEQ_START)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(186)
    defparam \DdrCtrl_CFG_SEQ_START~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_SEQ_START~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_CFG_SEQ_START~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_CFG_SEQ_START~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_CFG_SEQ_START~FF .SR_SYNC = 1'b0;
    defparam \DdrCtrl_CFG_SEQ_START~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_CFG_SEQ_START~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n92 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] ), 
           .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(186)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(150)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF  (.D(1'b1), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(150)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF  (.D(n162), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF  (.D(\U0_DDR_Reset/u_ddr_reset_sequencer/n91 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] ), 
           .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(186)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF  (.D(n1158), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF  (.D(n1156), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF  (.D(n1142), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF  (.D(n1140), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF  (.D(n1008), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF  (.D(n1006), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF  (.D(n989), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF  (.D(n971), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF  (.D(n969), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF  (.D(n967), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF  (.D(n965), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF  (.D(n963), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF  (.D(n961), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF  (.D(n959), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF  (.D(n957), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF  (.D(n955), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF  (.D(n953), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .SR_VALUE = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF  (.D(n951), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF  (.D(n950), .CE(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_CFG_RST_N), .Q(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(171)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .CLK_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .CE_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .SR_POLARITY = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .D_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .SR_SYNC = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .SR_VALUE = 1'b0;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/pCnt_value[0]~FF  (.D(\u_VsyHsyGenerator/pCnt_valueNext[0] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/pCnt_value[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/pCnt_value[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[0]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[0]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[0]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/frameCnt_value[0]~FF  (.D(\u_VsyHsyGenerator/frameCnt_valueNext[0] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/frameCnt_value[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/frameCnt_value[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[0]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[0]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[0]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/vsynDl[0]~FF  (.D(\u_VsyHsyGenerator/n402 ), 
           .CE(ceg_net2), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_VsyHsyGenerator/vsynDl[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/vsynDl[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/vsynDl[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/vsynDl[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/vsynDl[0]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/vsynDl[0]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/vsynDl[0]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/vsynDl[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/pCntInc~FF  (.D(\u_VsyHsyGenerator/when_MyTopLevel_l56 ), 
           .CE(ceg_net5), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_VsyHsyGenerator/pCntInc )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/pCntInc~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCntInc~FF .CE_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/pCntInc~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/pCntInc~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCntInc~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/pCntInc~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/pCntInc~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/hsynDl[0]~FF  (.D(\u_VsyHsyGenerator/n519 ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/hsynDl[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/hsynDl[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynDl[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynDl[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/hsynDl[0]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynDl[0]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/hsynDl[0]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/hsynDl[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/hsynCnt_value[0]~FF  (.D(\u_VsyHsyGenerator/hsynCnt_valueNext[0] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/hsynCnt_value[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/hsynCnt_value[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[0]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[0]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[0]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/pCnt_value[1]~FF  (.D(\u_VsyHsyGenerator/pCnt_valueNext[1] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/pCnt_value[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/pCnt_value[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[1]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[1]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[1]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/pCnt_value[2]~FF  (.D(\u_VsyHsyGenerator/pCnt_valueNext[2] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/pCnt_value[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/pCnt_value[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[2]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[2]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[2]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/pCnt_value[3]~FF  (.D(\u_VsyHsyGenerator/pCnt_valueNext[3] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/pCnt_value[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/pCnt_value[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[3]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[3]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[3]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/pCnt_value[4]~FF  (.D(\u_VsyHsyGenerator/pCnt_valueNext[4] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/pCnt_value[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/pCnt_value[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[4]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[4]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[4]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/pCnt_value[5]~FF  (.D(\u_VsyHsyGenerator/pCnt_valueNext[5] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/pCnt_value[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/pCnt_value[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[5]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[5]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[5]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/pCnt_value[6]~FF  (.D(\u_VsyHsyGenerator/pCnt_valueNext[6] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/pCnt_value[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/pCnt_value[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[6]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[6]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[6]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/pCnt_value[7]~FF  (.D(\u_VsyHsyGenerator/pCnt_valueNext[7] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/pCnt_value[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/pCnt_value[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[7]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[7]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[7]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/pCnt_value[8]~FF  (.D(\u_VsyHsyGenerator/pCnt_valueNext[8] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/pCnt_value[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/pCnt_value[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[8]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[8]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[8]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/pCnt_value[9]~FF  (.D(\u_VsyHsyGenerator/pCnt_valueNext[9] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/pCnt_value[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/pCnt_value[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[9]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[9]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[9]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/pCnt_value[10]~FF  (.D(\u_VsyHsyGenerator/pCnt_valueNext[10] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/pCnt_value[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/pCnt_value[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[10]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/pCnt_value[10]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[10]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/pCnt_value[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/frameCnt_value[1]~FF  (.D(\u_VsyHsyGenerator/frameCnt_valueNext[1] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/frameCnt_value[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/frameCnt_value[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[1]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[1]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[1]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/frameCnt_value[2]~FF  (.D(\u_VsyHsyGenerator/frameCnt_valueNext[2] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/frameCnt_value[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/frameCnt_value[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[2]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[2]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[2]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/frameCnt_value[3]~FF  (.D(\u_VsyHsyGenerator/frameCnt_valueNext[3] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/frameCnt_value[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/frameCnt_value[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[3]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[3]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[3]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/frameCnt_value[4]~FF  (.D(\u_VsyHsyGenerator/frameCnt_valueNext[4] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/frameCnt_value[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/frameCnt_value[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[4]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[4]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[4]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/frameCnt_value[5]~FF  (.D(\u_VsyHsyGenerator/frameCnt_valueNext[5] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/frameCnt_value[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/frameCnt_value[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[5]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[5]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[5]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/frameCnt_value[6]~FF  (.D(\u_VsyHsyGenerator/frameCnt_valueNext[6] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/frameCnt_value[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/frameCnt_value[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[6]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[6]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[6]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/frameCnt_value[7]~FF  (.D(\u_VsyHsyGenerator/frameCnt_valueNext[7] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/frameCnt_value[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/frameCnt_value[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[7]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[7]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[7]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/frameCnt_value[8]~FF  (.D(\u_VsyHsyGenerator/frameCnt_valueNext[8] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/frameCnt_value[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/frameCnt_value[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[8]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[8]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[8]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/frameCnt_value[9]~FF  (.D(\u_VsyHsyGenerator/frameCnt_valueNext[9] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/frameCnt_value[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/frameCnt_value[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[9]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/frameCnt_value[9]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[9]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/frameCnt_value[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/vsynDl[1]~FF  (.D(\u_VsyHsyGenerator/vsynDl[0] ), 
           .CE(\u_VsyHsyGenerator/n681 ), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_VsyHsyGenerator/vsynDl[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/vsynDl[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/vsynDl[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/vsynDl[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/vsynDl[1]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/vsynDl[1]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/vsynDl[1]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/vsynDl[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/vsynDl[2]~FF  (.D(\u_VsyHsyGenerator/vsynDl[1] ), 
           .CE(\u_VsyHsyGenerator/n681 ), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), 
           .Q(\u_VsyHsyGenerator/vsynDl[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/vsynDl[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/vsynDl[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/vsynDl[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/vsynDl[2]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/vsynDl[2]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/vsynDl[2]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/vsynDl[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XYCrop_frame_vsync~FF  (.D(\u_VsyHsyGenerator/vsynDl[2] ), .CE(\u_VsyHsyGenerator/n681 ), 
           .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(XYCrop_frame_vsync)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \XYCrop_frame_vsync~FF .CLK_POLARITY = 1'b1;
    defparam \XYCrop_frame_vsync~FF .CE_POLARITY = 1'b1;
    defparam \XYCrop_frame_vsync~FF .SR_POLARITY = 1'b0;
    defparam \XYCrop_frame_vsync~FF .D_POLARITY = 1'b1;
    defparam \XYCrop_frame_vsync~FF .SR_SYNC = 1'b0;
    defparam \XYCrop_frame_vsync~FF .SR_VALUE = 1'b0;
    defparam \XYCrop_frame_vsync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/hsynDl[1]~FF  (.D(\u_VsyHsyGenerator/n416 ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/hsynDl[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/hsynDl[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynDl[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynDl[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/hsynDl[1]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynDl[1]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/hsynDl[1]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/hsynDl[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/hsynDl[2]~FF  (.D(\u_VsyHsyGenerator/n415 ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/hsynDl[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/hsynDl[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynDl[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynDl[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/hsynDl[2]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynDl[2]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/hsynDl[2]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/hsynDl[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \XYCrop_frame_href~FF  (.D(\u_VsyHsyGenerator/n414 ), .CE(1'b1), 
           .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(XYCrop_frame_href)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \XYCrop_frame_href~FF .CLK_POLARITY = 1'b1;
    defparam \XYCrop_frame_href~FF .CE_POLARITY = 1'b1;
    defparam \XYCrop_frame_href~FF .SR_POLARITY = 1'b0;
    defparam \XYCrop_frame_href~FF .D_POLARITY = 1'b1;
    defparam \XYCrop_frame_href~FF .SR_SYNC = 1'b0;
    defparam \XYCrop_frame_href~FF .SR_VALUE = 1'b0;
    defparam \XYCrop_frame_href~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/hsynCnt_value[1]~FF  (.D(\u_VsyHsyGenerator/hsynCnt_valueNext[1] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/hsynCnt_value[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/hsynCnt_value[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[1]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[1]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[1]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/hsynCnt_value[2]~FF  (.D(\u_VsyHsyGenerator/hsynCnt_valueNext[2] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/hsynCnt_value[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/hsynCnt_value[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[2]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[2]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[2]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/hsynCnt_value[3]~FF  (.D(\u_VsyHsyGenerator/hsynCnt_valueNext[3] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/hsynCnt_value[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/hsynCnt_value[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[3]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[3]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[3]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/hsynCnt_value[4]~FF  (.D(\u_VsyHsyGenerator/hsynCnt_valueNext[4] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/hsynCnt_value[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/hsynCnt_value[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[4]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[4]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[4]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/hsynCnt_value[5]~FF  (.D(\u_VsyHsyGenerator/hsynCnt_valueNext[5] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/hsynCnt_value[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/hsynCnt_value[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[5]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[5]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[5]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/hsynCnt_value[6]~FF  (.D(\u_VsyHsyGenerator/hsynCnt_valueNext[6] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/hsynCnt_value[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/hsynCnt_value[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[6]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[6]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[6]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/hsynCnt_value[7]~FF  (.D(\u_VsyHsyGenerator/hsynCnt_valueNext[7] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/hsynCnt_value[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/hsynCnt_value[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[7]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[7]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[7]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/hsynCnt_value[8]~FF  (.D(\u_VsyHsyGenerator/hsynCnt_valueNext[8] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/hsynCnt_value[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/hsynCnt_value[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[8]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[8]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[8]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_VsyHsyGenerator/hsynCnt_value[9]~FF  (.D(\u_VsyHsyGenerator/hsynCnt_valueNext[9] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_VsyHsyGenerator/hsynCnt_value[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(246)
    defparam \u_VsyHsyGenerator/hsynCnt_value[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[9]~FF .D_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/hsynCnt_value[9]~FF .SR_SYNC = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[9]~FF .SR_VALUE = 1'b0;
    defparam \u_VsyHsyGenerator/hsynCnt_value[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wframe_vsync_dly[0]~FF  (.D(XYCrop_frame_vsync), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/wframe_vsync_dly[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(77)
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wframe_index[1]~FF  (.D(\u_axi4_ctrl/n323 ), .CE(\u_axi4_ctrl/equal_37/n3 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/wframe_index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(175)
    defparam \u_axi4_ctrl/wframe_index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_index[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_index[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_index[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_index[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wframe_index[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wframe_index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rframe_vsync_dly[0]~FF  (.D(\u_lcd_driver/n108 ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rframe_vsync_dly[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(77)
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wfifo_cnt[0]~FF  (.D(\u_axi4_ctrl/n96 ), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1476 ), .Q(\u_axi4_ctrl/wfifo_cnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(94)
    defparam \u_axi4_ctrl/wfifo_cnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[0]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wfifo_rst~FF  (.D(\u_axi4_ctrl/equal_28/n9 ), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/wfifo_rst )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(109)
    defparam \u_axi4_ctrl/wfifo_rst~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_rst~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_rst~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wfifo_rst~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_rst~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wfifo_rst~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/wfifo_rst~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wframe_index[0]~FF  (.D(\u_axi4_ctrl/n324 ), .CE(\u_axi4_ctrl/equal_37/n3 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/wframe_index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(175)
    defparam \u_axi4_ctrl/wframe_index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_index[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_index[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_index[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_index[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wframe_index[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wframe_index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rframe_index[0]~FF  (.D(\u_axi4_ctrl/n343 ), .CE(\u_axi4_ctrl/equal_46/n3 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rframe_index[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(195)
    defparam \u_axi4_ctrl/rframe_index[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_index[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_index[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rframe_index[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/state[0]~FF  (.D(\u_axi4_ctrl/n396 ), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/state[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(266)
    defparam \u_axi4_ctrl/state[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/state[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/state[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/state[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wframe_vsync_dly[1]~FF  (.D(\u_axi4_ctrl/wframe_vsync_dly[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/wframe_vsync_dly[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(77)
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_WSTRB_0[15]~FF  (.D(1'b1), .CE(1'b1), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(DdrCtrl_ABURST_0[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(59)
    defparam \DdrCtrl_WSTRB_0[15]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_WSTRB_0[15]~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_WSTRB_0[15]~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_WSTRB_0[15]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_WSTRB_0[15]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_WSTRB_0[15]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_WSTRB_0[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_ATYPE_0~FF  (.D(1'b1), .CE(\u_axi4_ctrl/n412 ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/n1483 ), .Q(DdrCtrl_ATYPE_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(281)
    defparam \DdrCtrl_ATYPE_0~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_ATYPE_0~FF .CE_POLARITY = 1'b1;
    defparam \DdrCtrl_ATYPE_0~FF .SR_POLARITY = 1'b1;
    defparam \DdrCtrl_ATYPE_0~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_ATYPE_0~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_ATYPE_0~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_ATYPE_0~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wframe_vsync_dly[3]~FF  (.D(\u_axi4_ctrl/wframe_vsync_dly[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/wframe_vsync_dly[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(77)
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/wfifo_rst ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(499)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/wfifo_rst ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(499)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/wfifo_rst ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(492)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wfifo_cnt[4]~FF  (.D(\u_axi4_ctrl/n92 ), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1476 ), .Q(\u_axi4_ctrl/wfifo_cnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(94)
    defparam \u_axi4_ctrl/wfifo_cnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[4]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wfifo_cnt[3]~FF  (.D(\u_axi4_ctrl/n93 ), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1476 ), .Q(\u_axi4_ctrl/wfifo_cnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(94)
    defparam \u_axi4_ctrl/wfifo_cnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[3]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[0]~FF  (.D(\u_axi4_ctrl/wdata_cnt_dly[0] ), 
           .CE(\u_axi4_ctrl/n370 ), .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), 
           .Q(\u_axi4_ctrl/wdata_cnt_dly[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(345)
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[1]~FF  (.D(\u_axi4_ctrl/n1551 ), .CE(\u_axi4_ctrl/n386 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(396)
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[0]~FF  (.D(\u_axi4_ctrl/rdata_cnt_dly[0] ), 
           .CE(\u_axi4_ctrl/n386 ), .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), 
           .Q(\u_axi4_ctrl/rdata_cnt_dly[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(396)
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wfifo_cnt[2]~FF  (.D(\u_axi4_ctrl/n94 ), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1476 ), .Q(\u_axi4_ctrl/wfifo_cnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(94)
    defparam \u_axi4_ctrl/wfifo_cnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[2]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wfifo_cnt[1]~FF  (.D(\u_axi4_ctrl/n95 ), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1476 ), .Q(\u_axi4_ctrl/wfifo_cnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(94)
    defparam \u_axi4_ctrl/wfifo_cnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/wfifo_cnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rframe_vsync_dly[3]~FF  (.D(\u_axi4_ctrl/rframe_vsync_dly[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rframe_vsync_dly[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(77)
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rframe_vsync_dly[2]~FF  (.D(\u_axi4_ctrl/rframe_vsync_dly[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rframe_vsync_dly[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(77)
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wenb~FF  (.D(\u_axi4_ctrl/n386 ), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rfifo_wenb )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(430)
    defparam \u_axi4_ctrl/rfifo_wenb~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wenb~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wenb~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wenb~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wenb~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wenb~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wenb~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rframe_vsync_dly[1]~FF  (.D(\u_axi4_ctrl/rframe_vsync_dly[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rframe_vsync_dly[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(77)
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rframe_vsync_dly[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[0]~FF  (.D(DdrCtrl_RDATA_0[0]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wframe_vsync_dly[2]~FF  (.D(\u_axi4_ctrl/wframe_vsync_dly[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/wframe_vsync_dly[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(77)
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wframe_vsync_dly[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF  (.D(n401), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF  (.D(n420), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\clk_12M_i~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF  (.D(n418), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wfifo_empty~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CE(ceg_net12), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/wfifo_empty )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1090)
    defparam \u_axi4_ctrl/wfifo_empty~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_empty~FF .CE_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wfifo_empty~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wfifo_empty~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wfifo_empty~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/wfifo_empty~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/wfifo_empty~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF  (.D(n380), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\clk_12M_i~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF  (.D(n422), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF  (.D(n381), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\clk_12M_i~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF  (.D(n397), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\clk_12M_i~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[0] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF  (.D(n405), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF  (.D(n409), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF  (.D(n413), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF  (.D(n415), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF  (.D(n569), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF  (.D(n597), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF  (.D(n344), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF  (.D(n342), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF  (.D(n340), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF  (.D(n338), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF  (.D(n336), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF  (.D(n334), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8]~FF  (.D(n332), .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[9]~FF  (.D(n331), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[9] ), 
           .CE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[1] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[8] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[8] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[9] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[10] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[11] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[2] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[0] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[1] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][0] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][1] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][2] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][12] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF  (.D(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0] ), 
           .CE(1'b1), .CLK(\clk_12M_i~O ), .SR(\u_axi4_ctrl/wfifo_rst ), 
           .Q(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(492)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(499)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(499)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF  (.D(1'b0), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(492)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_empty~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CE(ceg_net19), .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/rfifo_empty )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1090)
    defparam \u_axi4_ctrl/rfifo_empty~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_empty~FF .CE_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rfifo_empty~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_empty~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rfifo_empty~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/rfifo_empty~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/rfifo_empty~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\tx_slowclk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[0] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF  (.D(n747), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF  (.D(n754), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF  (.D(n295), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF  (.D(n293), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF  (.D(n291), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF  (.D(n289), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF  (.D(n287), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF  (.D(n286), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), .CLK(\Axi_Clk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1273)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF  (.D(n758), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF  (.D(n284), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF  (.D(n282), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF  (.D(n280), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF  (.D(n278), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF  (.D(n276), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF  (.D(n274), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF  (.D(n272), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF  (.D(n270), .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), 
           .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF  (.D(n268), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\tx_slowclk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[11]~FF  (.D(n267), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\tx_slowclk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\tx_slowclk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\tx_slowclk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\tx_slowclk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\tx_slowclk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\tx_slowclk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\tx_slowclk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\tx_slowclk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\tx_slowclk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[11] ), 
           .CE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .CLK(\tx_slowclk~O ), 
           .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1284)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1316)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[1] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1325)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[8] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[9] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[10] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[11] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.rd_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1339)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] ), 
           .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1351)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_r[11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][3] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][7] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][8] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][9] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][10] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.xrd2wr_addr_sync/pipe_reg[0][11] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[5] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[4] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[3] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[2] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[6] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[0] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[1] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[7] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_r[8] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][0] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][1] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][2] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][3] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][4] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][5] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][6] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][7] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.wr2rd_addr_sync/pipe_reg[0][8] ), 
           .CE(1'b1), .CLK(\tx_slowclk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(133)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF  (.D(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[0] ), 
           .CE(1'b1), .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0, async_reg="true" */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(492)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/genblk2.wr_rst[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rframe_index[1]~FF  (.D(\u_axi4_ctrl/n342 ), .CE(\u_axi4_ctrl/equal_46/n3 ), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/rframe_index[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(195)
    defparam \u_axi4_ctrl/rframe_index[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_index[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rframe_index[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[1]~FF .SR_VALUE = 1'b1;
    defparam \u_axi4_ctrl/rframe_index[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/state[1]~FF  (.D(\u_axi4_ctrl/n1616 ), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1623 ), .Q(\u_axi4_ctrl/state[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(266)
    defparam \u_axi4_ctrl/state[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/state[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/state[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/state[2]~FF  (.D(\u_axi4_ctrl/n394 ), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_axi4_ctrl/state[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(266)
    defparam \u_axi4_ctrl/state[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/state[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/state[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/state[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/state[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[10]~FF  (.D(\u_axi4_ctrl/awaddr[10] ), .CE(\u_axi4_ctrl/n376 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1476 ), .Q(\u_axi4_ctrl/awaddr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl/awaddr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[10]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/awaddr[10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[11]~FF  (.D(n411), .CE(\u_axi4_ctrl/n376 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1476 ), .Q(\u_axi4_ctrl/awaddr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl/awaddr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[12]~FF  (.D(n721), .CE(\u_axi4_ctrl/n376 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1476 ), .Q(\u_axi4_ctrl/awaddr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl/awaddr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[13]~FF  (.D(n719), .CE(\u_axi4_ctrl/n376 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1476 ), .Q(\u_axi4_ctrl/awaddr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl/awaddr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[13]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[13]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[13]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[14]~FF  (.D(n717), .CE(\u_axi4_ctrl/n376 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1476 ), .Q(\u_axi4_ctrl/awaddr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl/awaddr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[14]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[14]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[14]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[15]~FF  (.D(n715), .CE(\u_axi4_ctrl/n376 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1476 ), .Q(\u_axi4_ctrl/awaddr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl/awaddr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[15]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[15]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[15]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[16]~FF  (.D(n713), .CE(\u_axi4_ctrl/n376 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1476 ), .Q(\u_axi4_ctrl/awaddr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl/awaddr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[16]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[16]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[16]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[17]~FF  (.D(n593), .CE(\u_axi4_ctrl/n376 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1476 ), .Q(\u_axi4_ctrl/awaddr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl/awaddr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[17]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[17]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[17]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[18]~FF  (.D(n565), .CE(\u_axi4_ctrl/n376 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1476 ), .Q(\u_axi4_ctrl/awaddr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl/awaddr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[18]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[18]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[18]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[19]~FF  (.D(n563), .CE(\u_axi4_ctrl/n376 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1476 ), .Q(\u_axi4_ctrl/awaddr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl/awaddr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[19]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[19]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[19]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[20]~FF  (.D(n559), .CE(\u_axi4_ctrl/n376 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1476 ), .Q(\u_axi4_ctrl/awaddr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl/awaddr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[20]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[20]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[20]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[21]~FF  (.D(n554), .CE(\u_axi4_ctrl/n376 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1476 ), .Q(\u_axi4_ctrl/awaddr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl/awaddr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[21]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[21]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[21]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[22]~FF  (.D(n552), .CE(\u_axi4_ctrl/n376 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1476 ), .Q(\u_axi4_ctrl/awaddr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl/awaddr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[22]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[22]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[22]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[22]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/awaddr[23]~FF  (.D(n551), .CE(\u_axi4_ctrl/n376 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1476 ), .Q(\u_axi4_ctrl/awaddr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(298)
    defparam \u_axi4_ctrl/awaddr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[23]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[23]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/awaddr[23]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/awaddr[23]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/awaddr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[10]~FF  (.D(\u_axi4_ctrl/araddr[10] ), .CE(\u_axi4_ctrl/n388 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1485 ), .Q(\u_axi4_ctrl/araddr[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/araddr[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[10]~FF .D_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/araddr[10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[11]~FF  (.D(n460), .CE(\u_axi4_ctrl/n388 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1485 ), .Q(\u_axi4_ctrl/araddr[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/araddr[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[12]~FF  (.D(n470), .CE(\u_axi4_ctrl/n388 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1485 ), .Q(\u_axi4_ctrl/araddr[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/araddr[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[13]~FF  (.D(n543), .CE(\u_axi4_ctrl/n388 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1485 ), .Q(\u_axi4_ctrl/araddr[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/araddr[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[13]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[13]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[13]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[14]~FF  (.D(n541), .CE(\u_axi4_ctrl/n388 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1485 ), .Q(\u_axi4_ctrl/araddr[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/araddr[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[14]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[14]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[14]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[15]~FF  (.D(n539), .CE(\u_axi4_ctrl/n388 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1485 ), .Q(\u_axi4_ctrl/araddr[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/araddr[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[15]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[15]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[15]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[16]~FF  (.D(n490), .CE(\u_axi4_ctrl/n388 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1485 ), .Q(\u_axi4_ctrl/araddr[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/araddr[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[16]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[16]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[16]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[17]~FF  (.D(n488), .CE(\u_axi4_ctrl/n388 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1485 ), .Q(\u_axi4_ctrl/araddr[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/araddr[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[17]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[17]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[17]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[18]~FF  (.D(n486), .CE(\u_axi4_ctrl/n388 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1485 ), .Q(\u_axi4_ctrl/araddr[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/araddr[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[18]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[18]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[18]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[19]~FF  (.D(n484), .CE(\u_axi4_ctrl/n388 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1485 ), .Q(\u_axi4_ctrl/araddr[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/araddr[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[19]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[19]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[19]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[20]~FF  (.D(n482), .CE(\u_axi4_ctrl/n388 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1485 ), .Q(\u_axi4_ctrl/araddr[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/araddr[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[20]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[20]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[20]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[21]~FF  (.D(n480), .CE(\u_axi4_ctrl/n388 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1485 ), .Q(\u_axi4_ctrl/araddr[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/araddr[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[21]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[21]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[21]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[22]~FF  (.D(n426), .CE(\u_axi4_ctrl/n388 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1485 ), .Q(\u_axi4_ctrl/araddr[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/araddr[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[22]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[22]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[22]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[22]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/araddr[23]~FF  (.D(n425), .CE(\u_axi4_ctrl/n388 ), 
           .CLK(\Axi_Clk~O ), .SR(\u_axi4_ctrl/n1485 ), .Q(\u_axi4_ctrl/araddr[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(315)
    defparam \u_axi4_ctrl/araddr[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[23]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[23]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/araddr[23]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/araddr[23]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/araddr[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[10]~FF  (.D(\u_axi4_ctrl/n704 ), .CE(ceg_net124), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(330)
    defparam \DdrCtrl_AADDR_0[10]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[10]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[10]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[10]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[10]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[10]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[11]~FF  (.D(\u_axi4_ctrl/n703 ), .CE(ceg_net124), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(330)
    defparam \DdrCtrl_AADDR_0[11]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[11]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[11]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[11]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[11]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[11]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[12]~FF  (.D(\u_axi4_ctrl/n702 ), .CE(ceg_net124), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(330)
    defparam \DdrCtrl_AADDR_0[12]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[12]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[12]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[12]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[12]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[12]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[13]~FF  (.D(\u_axi4_ctrl/n701 ), .CE(ceg_net124), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(330)
    defparam \DdrCtrl_AADDR_0[13]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[13]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[13]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[13]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[13]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[13]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[14]~FF  (.D(\u_axi4_ctrl/n700 ), .CE(ceg_net124), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(330)
    defparam \DdrCtrl_AADDR_0[14]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[14]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[14]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[14]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[14]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[14]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[15]~FF  (.D(\u_axi4_ctrl/n699 ), .CE(ceg_net124), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(330)
    defparam \DdrCtrl_AADDR_0[15]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[15]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[15]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[15]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[15]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[15]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[16]~FF  (.D(\u_axi4_ctrl/n698 ), .CE(ceg_net124), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(330)
    defparam \DdrCtrl_AADDR_0[16]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[16]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[16]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[16]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[16]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[16]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[17]~FF  (.D(\u_axi4_ctrl/n697 ), .CE(ceg_net124), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(330)
    defparam \DdrCtrl_AADDR_0[17]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[17]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[17]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[17]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[17]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[17]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[18]~FF  (.D(\u_axi4_ctrl/n696 ), .CE(ceg_net124), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(330)
    defparam \DdrCtrl_AADDR_0[18]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[18]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[18]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[18]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[18]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[18]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[19]~FF  (.D(\u_axi4_ctrl/n695 ), .CE(ceg_net124), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(330)
    defparam \DdrCtrl_AADDR_0[19]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[19]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[19]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[19]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[19]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[19]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[20]~FF  (.D(\u_axi4_ctrl/n694 ), .CE(ceg_net124), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(330)
    defparam \DdrCtrl_AADDR_0[20]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[20]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[20]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[20]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[20]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[20]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[21]~FF  (.D(\u_axi4_ctrl/n693 ), .CE(ceg_net124), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(330)
    defparam \DdrCtrl_AADDR_0[21]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[21]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[21]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[21]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[21]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[21]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[22]~FF  (.D(\u_axi4_ctrl/n692 ), .CE(ceg_net124), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(330)
    defparam \DdrCtrl_AADDR_0[22]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[22]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[22]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[22]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[22]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[22]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[23]~FF  (.D(\u_axi4_ctrl/n691 ), .CE(ceg_net124), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(330)
    defparam \DdrCtrl_AADDR_0[23]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[23]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[23]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[23]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[23]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[23]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[24]~FF  (.D(\u_axi4_ctrl/n690 ), .CE(ceg_net124), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(330)
    defparam \DdrCtrl_AADDR_0[24]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[24]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[24]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[24]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[24]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[24]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \DdrCtrl_AADDR_0[25]~FF  (.D(\u_axi4_ctrl/n689 ), .CE(ceg_net124), 
           .CLK(\Axi_Clk~O ), .SR(\Axi0ResetReg[2] ), .Q(DdrCtrl_AADDR_0[25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(330)
    defparam \DdrCtrl_AADDR_0[25]~FF .CLK_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[25]~FF .CE_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[25]~FF .SR_POLARITY = 1'b0;
    defparam \DdrCtrl_AADDR_0[25]~FF .D_POLARITY = 1'b1;
    defparam \DdrCtrl_AADDR_0[25]~FF .SR_SYNC = 1'b1;
    defparam \DdrCtrl_AADDR_0[25]~FF .SR_VALUE = 1'b0;
    defparam \DdrCtrl_AADDR_0[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[1]~FF  (.D(\u_axi4_ctrl/n1506 ), .CE(\u_axi4_ctrl/n370 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(345)
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[2]~FF  (.D(\u_axi4_ctrl/n1511 ), .CE(\u_axi4_ctrl/n370 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(345)
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[3]~FF  (.D(\u_axi4_ctrl/n1516 ), .CE(\u_axi4_ctrl/n370 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(345)
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[4]~FF  (.D(\u_axi4_ctrl/n1521 ), .CE(\u_axi4_ctrl/n370 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(345)
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[5]~FF  (.D(\u_axi4_ctrl/n1526 ), .CE(\u_axi4_ctrl/n370 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(345)
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[6]~FF  (.D(\u_axi4_ctrl/n1531 ), .CE(\u_axi4_ctrl/n370 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(345)
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[7]~FF  (.D(\u_axi4_ctrl/n1536 ), .CE(\u_axi4_ctrl/n370 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(345)
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/wdata_cnt_dly[8]~FF  (.D(\u_axi4_ctrl/n1541 ), .CE(\u_axi4_ctrl/n370 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_WVALID_0), .Q(\u_axi4_ctrl/wdata_cnt_dly[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(345)
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/wdata_cnt_dly[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[2]~FF  (.D(\u_axi4_ctrl/n1556 ), .CE(\u_axi4_ctrl/n386 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(396)
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[3]~FF  (.D(\u_axi4_ctrl/n1561 ), .CE(\u_axi4_ctrl/n386 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(396)
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[4]~FF  (.D(\u_axi4_ctrl/n1566 ), .CE(\u_axi4_ctrl/n386 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(396)
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[5]~FF  (.D(\u_axi4_ctrl/n1571 ), .CE(\u_axi4_ctrl/n386 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(396)
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[6]~FF  (.D(\u_axi4_ctrl/n1576 ), .CE(\u_axi4_ctrl/n386 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(396)
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[7]~FF  (.D(\u_axi4_ctrl/n1581 ), .CE(\u_axi4_ctrl/n386 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(396)
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rdata_cnt_dly[8]~FF  (.D(\u_axi4_ctrl/n1586 ), .CE(\u_axi4_ctrl/n386 ), 
           .CLK(\Axi_Clk~O ), .SR(DdrCtrl_RREADY_0), .Q(\u_axi4_ctrl/rdata_cnt_dly[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(396)
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rdata_cnt_dly[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[1]~FF  (.D(DdrCtrl_RDATA_0[1]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[2]~FF  (.D(DdrCtrl_RDATA_0[2]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[3]~FF  (.D(DdrCtrl_RDATA_0[3]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[4]~FF  (.D(DdrCtrl_RDATA_0[4]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[5]~FF  (.D(DdrCtrl_RDATA_0[5]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[6]~FF  (.D(DdrCtrl_RDATA_0[6]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[7]~FF  (.D(DdrCtrl_RDATA_0[7]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[8]~FF  (.D(DdrCtrl_RDATA_0[8]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[9]~FF  (.D(DdrCtrl_RDATA_0[9]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[10]~FF  (.D(DdrCtrl_RDATA_0[10]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[11]~FF  (.D(DdrCtrl_RDATA_0[11]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[12]~FF  (.D(DdrCtrl_RDATA_0[12]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[13]~FF  (.D(DdrCtrl_RDATA_0[13]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[14]~FF  (.D(DdrCtrl_RDATA_0[14]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[15]~FF  (.D(DdrCtrl_RDATA_0[15]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[16]~FF  (.D(DdrCtrl_RDATA_0[16]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[17]~FF  (.D(DdrCtrl_RDATA_0[17]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[18]~FF  (.D(DdrCtrl_RDATA_0[18]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[19]~FF  (.D(DdrCtrl_RDATA_0[19]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[20]~FF  (.D(DdrCtrl_RDATA_0[20]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[21]~FF  (.D(DdrCtrl_RDATA_0[21]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[22]~FF  (.D(DdrCtrl_RDATA_0[22]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[23]~FF  (.D(DdrCtrl_RDATA_0[23]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[24]~FF  (.D(DdrCtrl_RDATA_0[24]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[25]~FF  (.D(DdrCtrl_RDATA_0[25]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[26]~FF  (.D(DdrCtrl_RDATA_0[26]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[27]~FF  (.D(DdrCtrl_RDATA_0[27]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[28]~FF  (.D(DdrCtrl_RDATA_0[28]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[29]~FF  (.D(DdrCtrl_RDATA_0[29]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[30]~FF  (.D(DdrCtrl_RDATA_0[30]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[31]~FF  (.D(DdrCtrl_RDATA_0[31]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[32]~FF  (.D(DdrCtrl_RDATA_0[32]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[33]~FF  (.D(DdrCtrl_RDATA_0[33]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[34]~FF  (.D(DdrCtrl_RDATA_0[34]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[35]~FF  (.D(DdrCtrl_RDATA_0[35]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[36]~FF  (.D(DdrCtrl_RDATA_0[36]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[37]~FF  (.D(DdrCtrl_RDATA_0[37]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[38]~FF  (.D(DdrCtrl_RDATA_0[38]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[39]~FF  (.D(DdrCtrl_RDATA_0[39]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[40]~FF  (.D(DdrCtrl_RDATA_0[40]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[41]~FF  (.D(DdrCtrl_RDATA_0[41]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[42]~FF  (.D(DdrCtrl_RDATA_0[42]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[43]~FF  (.D(DdrCtrl_RDATA_0[43]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[44]~FF  (.D(DdrCtrl_RDATA_0[44]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[45]~FF  (.D(DdrCtrl_RDATA_0[45]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[46]~FF  (.D(DdrCtrl_RDATA_0[46]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[47]~FF  (.D(DdrCtrl_RDATA_0[47]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[48]~FF  (.D(DdrCtrl_RDATA_0[48]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[49]~FF  (.D(DdrCtrl_RDATA_0[49]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[50]~FF  (.D(DdrCtrl_RDATA_0[50]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[51]~FF  (.D(DdrCtrl_RDATA_0[51]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[52]~FF  (.D(DdrCtrl_RDATA_0[52]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[53]~FF  (.D(DdrCtrl_RDATA_0[53]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[54]~FF  (.D(DdrCtrl_RDATA_0[54]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[55]~FF  (.D(DdrCtrl_RDATA_0[55]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[56]~FF  (.D(DdrCtrl_RDATA_0[56]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[57]~FF  (.D(DdrCtrl_RDATA_0[57]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[58]~FF  (.D(DdrCtrl_RDATA_0[58]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[59]~FF  (.D(DdrCtrl_RDATA_0[59]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[60]~FF  (.D(DdrCtrl_RDATA_0[60]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[61]~FF  (.D(DdrCtrl_RDATA_0[61]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[62]~FF  (.D(DdrCtrl_RDATA_0[62]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[63]~FF  (.D(DdrCtrl_RDATA_0[63]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[64]~FF  (.D(DdrCtrl_RDATA_0[64]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[65]~FF  (.D(DdrCtrl_RDATA_0[65]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[66]~FF  (.D(DdrCtrl_RDATA_0[66]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[67]~FF  (.D(DdrCtrl_RDATA_0[67]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[68]~FF  (.D(DdrCtrl_RDATA_0[68]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[69]~FF  (.D(DdrCtrl_RDATA_0[69]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[70]~FF  (.D(DdrCtrl_RDATA_0[70]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[71]~FF  (.D(DdrCtrl_RDATA_0[71]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[72]~FF  (.D(DdrCtrl_RDATA_0[72]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[73]~FF  (.D(DdrCtrl_RDATA_0[73]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[74]~FF  (.D(DdrCtrl_RDATA_0[74]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[75]~FF  (.D(DdrCtrl_RDATA_0[75]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[76]~FF  (.D(DdrCtrl_RDATA_0[76]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[77]~FF  (.D(DdrCtrl_RDATA_0[77]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[78]~FF  (.D(DdrCtrl_RDATA_0[78]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[79]~FF  (.D(DdrCtrl_RDATA_0[79]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[80]~FF  (.D(DdrCtrl_RDATA_0[80]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[81]~FF  (.D(DdrCtrl_RDATA_0[81]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[82]~FF  (.D(DdrCtrl_RDATA_0[82]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[82] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[83]~FF  (.D(DdrCtrl_RDATA_0[83]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[83] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[84]~FF  (.D(DdrCtrl_RDATA_0[84]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[84] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[85]~FF  (.D(DdrCtrl_RDATA_0[85]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[85] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[86]~FF  (.D(DdrCtrl_RDATA_0[86]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[86] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[87]~FF  (.D(DdrCtrl_RDATA_0[87]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[87] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[88]~FF  (.D(DdrCtrl_RDATA_0[88]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[88] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[89]~FF  (.D(DdrCtrl_RDATA_0[89]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[89] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[90]~FF  (.D(DdrCtrl_RDATA_0[90]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[90] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[91]~FF  (.D(DdrCtrl_RDATA_0[91]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[91] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[92]~FF  (.D(DdrCtrl_RDATA_0[92]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[92] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[93]~FF  (.D(DdrCtrl_RDATA_0[93]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[93] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[94]~FF  (.D(DdrCtrl_RDATA_0[94]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[94] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[95]~FF  (.D(DdrCtrl_RDATA_0[95]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[95] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[96]~FF  (.D(DdrCtrl_RDATA_0[96]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[96] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[97]~FF  (.D(DdrCtrl_RDATA_0[97]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[97] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[98]~FF  (.D(DdrCtrl_RDATA_0[98]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[98] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[99]~FF  (.D(DdrCtrl_RDATA_0[99]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[99] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[100]~FF  (.D(DdrCtrl_RDATA_0[100]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[100] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[101]~FF  (.D(DdrCtrl_RDATA_0[101]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[101] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[102]~FF  (.D(DdrCtrl_RDATA_0[102]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[102] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[103]~FF  (.D(DdrCtrl_RDATA_0[103]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[103] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[104]~FF  (.D(DdrCtrl_RDATA_0[104]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[104] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[105]~FF  (.D(DdrCtrl_RDATA_0[105]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[105] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[106]~FF  (.D(DdrCtrl_RDATA_0[106]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[106] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[107]~FF  (.D(DdrCtrl_RDATA_0[107]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[107] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[108]~FF  (.D(DdrCtrl_RDATA_0[108]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[108] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[109]~FF  (.D(DdrCtrl_RDATA_0[109]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[109] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[110]~FF  (.D(DdrCtrl_RDATA_0[110]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[110] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[111]~FF  (.D(DdrCtrl_RDATA_0[111]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[111] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[112]~FF  (.D(DdrCtrl_RDATA_0[112]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[112] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[113]~FF  (.D(DdrCtrl_RDATA_0[113]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[113] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[114]~FF  (.D(DdrCtrl_RDATA_0[114]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[114] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[115]~FF  (.D(DdrCtrl_RDATA_0[115]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[115] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[116]~FF  (.D(DdrCtrl_RDATA_0[116]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[116] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[117]~FF  (.D(DdrCtrl_RDATA_0[117]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[117] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[118]~FF  (.D(DdrCtrl_RDATA_0[118]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[118] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[119]~FF  (.D(DdrCtrl_RDATA_0[119]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[119] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[120]~FF  (.D(DdrCtrl_RDATA_0[120]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[120] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[120]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[121]~FF  (.D(DdrCtrl_RDATA_0[121]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[121] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[121]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[122]~FF  (.D(DdrCtrl_RDATA_0[122]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[122] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[122]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[123]~FF  (.D(DdrCtrl_RDATA_0[123]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[123] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[123]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[124]~FF  (.D(DdrCtrl_RDATA_0[124]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[124] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[124]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[125]~FF  (.D(DdrCtrl_RDATA_0[125]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[125] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[125]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[126]~FF  (.D(DdrCtrl_RDATA_0[126]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[126] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[126]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_axi4_ctrl/rfifo_wdata[127]~FF  (.D(DdrCtrl_RDATA_0[127]), .CE(1'b1), 
           .CLK(\Axi_Clk~O ), .SR(1'b0), .Q(\u_axi4_ctrl/rfifo_wdata[127] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(435)
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .CLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .CE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .SR_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .D_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .SR_SYNC = 1'b1;
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .SR_VALUE = 1'b0;
    defparam \u_axi4_ctrl/rfifo_wdata[127]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[0]~FF  (.D(\u_lcd_driver/n81 ), .CE(\u_lcd_driver/equal_15/n23 ), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/vcnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(92)
    defparam \u_lcd_driver/vcnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[0]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[0]~FF  (.D(\u_lcd_driver/n34 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/hcnt[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(75)
    defparam \u_lcd_driver/hcnt[0]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[0]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[0]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[0]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[0]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[0]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[1]~FF  (.D(\u_lcd_driver/n80 ), .CE(\u_lcd_driver/equal_15/n23 ), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/vcnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(92)
    defparam \u_lcd_driver/vcnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[1]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[2]~FF  (.D(\u_lcd_driver/n79 ), .CE(\u_lcd_driver/equal_15/n23 ), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/vcnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(92)
    defparam \u_lcd_driver/vcnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[2]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[3]~FF  (.D(\u_lcd_driver/n78 ), .CE(\u_lcd_driver/equal_15/n23 ), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/vcnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(92)
    defparam \u_lcd_driver/vcnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[3]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[4]~FF  (.D(\u_lcd_driver/n77 ), .CE(\u_lcd_driver/equal_15/n23 ), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/vcnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(92)
    defparam \u_lcd_driver/vcnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[4]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[5]~FF  (.D(\u_lcd_driver/n76 ), .CE(\u_lcd_driver/equal_15/n23 ), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/vcnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(92)
    defparam \u_lcd_driver/vcnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[5]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[6]~FF  (.D(\u_lcd_driver/n75 ), .CE(\u_lcd_driver/equal_15/n23 ), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/vcnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(92)
    defparam \u_lcd_driver/vcnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[6]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[7]~FF  (.D(\u_lcd_driver/n74 ), .CE(\u_lcd_driver/equal_15/n23 ), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/vcnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(92)
    defparam \u_lcd_driver/vcnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[7]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[8]~FF  (.D(\u_lcd_driver/n73 ), .CE(\u_lcd_driver/equal_15/n23 ), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/vcnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(92)
    defparam \u_lcd_driver/vcnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[8]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[9]~FF  (.D(\u_lcd_driver/n72 ), .CE(\u_lcd_driver/equal_15/n23 ), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/vcnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(92)
    defparam \u_lcd_driver/vcnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[9]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[10]~FF  (.D(\u_lcd_driver/n71 ), .CE(\u_lcd_driver/equal_15/n23 ), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/vcnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(92)
    defparam \u_lcd_driver/vcnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[10]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/vcnt[11]~FF  (.D(\u_lcd_driver/n70 ), .CE(\u_lcd_driver/equal_15/n23 ), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/vcnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(92)
    defparam \u_lcd_driver/vcnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[11]~FF .CE_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/vcnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/vcnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/vcnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/vcnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[1]~FF  (.D(\u_lcd_driver/n33 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/hcnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(75)
    defparam \u_lcd_driver/hcnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[1]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[1]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[1]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[1]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[2]~FF  (.D(\u_lcd_driver/n32 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/hcnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(75)
    defparam \u_lcd_driver/hcnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[2]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[2]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[2]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[2]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[3]~FF  (.D(\u_lcd_driver/n31 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/hcnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(75)
    defparam \u_lcd_driver/hcnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[3]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[3]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[3]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[3]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[4]~FF  (.D(\u_lcd_driver/n30 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/hcnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(75)
    defparam \u_lcd_driver/hcnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[4]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[4]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[4]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[4]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[5]~FF  (.D(\u_lcd_driver/n29 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/hcnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(75)
    defparam \u_lcd_driver/hcnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[5]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[5]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[5]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[5]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[6]~FF  (.D(\u_lcd_driver/n28 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/hcnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(75)
    defparam \u_lcd_driver/hcnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[6]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[6]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[6]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[6]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[7]~FF  (.D(\u_lcd_driver/n27 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/hcnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(75)
    defparam \u_lcd_driver/hcnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[7]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[7]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[7]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[7]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[8]~FF  (.D(\u_lcd_driver/n26 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/hcnt[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(75)
    defparam \u_lcd_driver/hcnt[8]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[8]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[8]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[8]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[8]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[8]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[9]~FF  (.D(\u_lcd_driver/n25 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/hcnt[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(75)
    defparam \u_lcd_driver/hcnt[9]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[9]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[9]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[9]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[9]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[9]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[10]~FF  (.D(\u_lcd_driver/n24 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/hcnt[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(75)
    defparam \u_lcd_driver/hcnt[10]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[10]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[10]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[10]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[10]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[10]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \u_lcd_driver/hcnt[11]~FF  (.D(\u_lcd_driver/n23 ), .CE(1'b1), 
           .CLK(\tx_slowclk~O ), .SR(\Axi0ResetReg[2] ), .Q(\u_lcd_driver/hcnt[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(75)
    defparam \u_lcd_driver/hcnt[11]~FF .CLK_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[11]~FF .CE_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[11]~FF .SR_POLARITY = 1'b0;
    defparam \u_lcd_driver/hcnt[11]~FF .D_POLARITY = 1'b1;
    defparam \u_lcd_driver/hcnt[11]~FF .SR_SYNC = 1'b0;
    defparam \u_lcd_driver/hcnt[11]~FF .SR_VALUE = 1'b0;
    defparam \u_lcd_driver/hcnt[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[1]~FF  (.D(n1171), .CE(n6_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(99)
    defparam \PowerOnResetCnt[1]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[1]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[2]~FF  (.D(n1169), .CE(n6_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(99)
    defparam \PowerOnResetCnt[2]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[2]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[3]~FF  (.D(n1167), .CE(n6_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(99)
    defparam \PowerOnResetCnt[3]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[3]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[4]~FF  (.D(n1165), .CE(n6_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(99)
    defparam \PowerOnResetCnt[4]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[4]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[5]~FF  (.D(n1163), .CE(n6_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(99)
    defparam \PowerOnResetCnt[5]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[5]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[6]~FF  (.D(n1161), .CE(n6_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(99)
    defparam \PowerOnResetCnt[6]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[6]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \PowerOnResetCnt[7]~FF  (.D(n1160), .CE(n6_2), .CLK(\Axi_Clk~O ), 
           .SR(1'b0), .Q(\PowerOnResetCnt[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(99)
    defparam \PowerOnResetCnt[7]~FF .CLK_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .CE_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .SR_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .D_POLARITY = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .SR_SYNC = 1'b1;
    defparam \PowerOnResetCnt[7]~FF .SR_VALUE = 1'b0;
    defparam \PowerOnResetCnt[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0] ), 
            .I1(1'b0), .CI(n2552), .O(n162), .CO(n163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_24/i1  (.I0(\u_VsyHsyGenerator/hsynCnt_value[0] ), 
            .I1(n1405), .CI(1'b0), .O(n176), .CO(n177)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(102)
    defparam \u_VsyHsyGenerator/add_24/i1 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_24/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_31/i1  (.I0(\u_VsyHsyGenerator/pCnt_value[0] ), 
            .I1(\u_VsyHsyGenerator/pCntInc ), .CI(1'b0), .O(n198), .CO(n199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(129)
    defparam \u_VsyHsyGenerator/add_31/i1 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_31/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_39/i1  (.I0(\u_VsyHsyGenerator/frameCnt_value[0] ), 
            .I1(n1429), .CI(1'b0), .O(n200), .CO(n201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(158)
    defparam \u_VsyHsyGenerator/add_39/i1 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_39/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_17/i12  (.I0(\u_lcd_driver/vcnt[11] ), .I1(1'b0), 
            .CI(n218), .O(n216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(89)
    defparam \u_lcd_driver/add_17/i12 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_17/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_17/i11  (.I0(\u_lcd_driver/vcnt[10] ), .I1(1'b0), 
            .CI(n220), .O(n217), .CO(n218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(89)
    defparam \u_lcd_driver/add_17/i11 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_17/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_17/i10  (.I0(\u_lcd_driver/vcnt[9] ), .I1(1'b0), 
            .CI(n222), .O(n219), .CO(n220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(89)
    defparam \u_lcd_driver/add_17/i10 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_17/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_17/i9  (.I0(\u_lcd_driver/vcnt[8] ), .I1(1'b0), 
            .CI(n224), .O(n221), .CO(n222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(89)
    defparam \u_lcd_driver/add_17/i9 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_17/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_17/i8  (.I0(\u_lcd_driver/vcnt[7] ), .I1(1'b0), 
            .CI(n226), .O(n223), .CO(n224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(89)
    defparam \u_lcd_driver/add_17/i8 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_17/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_17/i7  (.I0(\u_lcd_driver/vcnt[6] ), .I1(1'b0), 
            .CI(n228), .O(n225), .CO(n226)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(89)
    defparam \u_lcd_driver/add_17/i7 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_17/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_17/i6  (.I0(\u_lcd_driver/vcnt[5] ), .I1(1'b0), 
            .CI(n230), .O(n227), .CO(n228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(89)
    defparam \u_lcd_driver/add_17/i6 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_17/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_17/i5  (.I0(\u_lcd_driver/vcnt[4] ), .I1(1'b0), 
            .CI(n232), .O(n229), .CO(n230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(89)
    defparam \u_lcd_driver/add_17/i5 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_17/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_17/i4  (.I0(\u_lcd_driver/vcnt[3] ), .I1(1'b0), 
            .CI(n234), .O(n231), .CO(n232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(89)
    defparam \u_lcd_driver/add_17/i4 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_17/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_17/i3  (.I0(\u_lcd_driver/vcnt[2] ), .I1(1'b0), 
            .CI(n1138), .O(n233), .CO(n234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(89)
    defparam \u_lcd_driver/add_17/i3 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_17/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i12  (.I0(\u_lcd_driver/hcnt[11] ), .I1(1'b0), 
            .CI(n237), .O(n235)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(72)
    defparam \u_lcd_driver/add_7/i12 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i11  (.I0(\u_lcd_driver/hcnt[10] ), .I1(1'b0), 
            .CI(n239), .O(n236), .CO(n237)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(72)
    defparam \u_lcd_driver/add_7/i11 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i10  (.I0(\u_lcd_driver/hcnt[9] ), .I1(1'b0), 
            .CI(n241), .O(n238), .CO(n239)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(72)
    defparam \u_lcd_driver/add_7/i10 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i9  (.I0(\u_lcd_driver/hcnt[8] ), .I1(1'b0), 
            .CI(n243), .O(n240), .CO(n241)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(72)
    defparam \u_lcd_driver/add_7/i9 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i8  (.I0(\u_lcd_driver/hcnt[7] ), .I1(1'b0), 
            .CI(n245), .O(n242), .CO(n243)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(72)
    defparam \u_lcd_driver/add_7/i8 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i7  (.I0(\u_lcd_driver/hcnt[6] ), .I1(1'b0), 
            .CI(n247), .O(n244), .CO(n245)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(72)
    defparam \u_lcd_driver/add_7/i7 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i6  (.I0(\u_lcd_driver/hcnt[5] ), .I1(1'b0), 
            .CI(n249), .O(n246), .CO(n247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(72)
    defparam \u_lcd_driver/add_7/i6 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i5  (.I0(\u_lcd_driver/hcnt[4] ), .I1(1'b0), 
            .CI(n251), .O(n248), .CO(n249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(72)
    defparam \u_lcd_driver/add_7/i5 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i4  (.I0(\u_lcd_driver/hcnt[3] ), .I1(1'b0), 
            .CI(n253), .O(n250), .CO(n251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(72)
    defparam \u_lcd_driver/add_7/i4 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i3  (.I0(\u_lcd_driver/hcnt[2] ), .I1(1'b0), 
            .CI(n777), .O(n252), .CO(n253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(72)
    defparam \u_lcd_driver/add_7/i3 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i8  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10] ), 
            .CI(n256), .O(n254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i7  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9] ), 
            .CI(n258), .O(n255), .CO(n256)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i6  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] ), 
            .CI(n260), .O(n257), .CO(n258)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i5  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] ), 
            .CI(n262), .O(n259), .CO(n260)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i4  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] ), 
            .CI(n264), .O(n261), .CO(n262)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i3  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] ), 
            .CI(n266), .O(n263), .CO(n264)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i2  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] ), 
            .CI(n762), .O(n265), .CO(n266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i12  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[11] ), 
            .I1(1'b0), .CI(n269), .O(n267)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i12 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i11  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] ), 
            .I1(1'b0), .CI(n271), .O(n268), .CO(n269)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i11 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i10  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] ), 
            .I1(1'b0), .CI(n273), .O(n270), .CO(n271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i10 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i9  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] ), 
            .I1(1'b0), .CI(n275), .O(n272), .CO(n273)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i8  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] ), 
            .I1(1'b0), .CI(n277), .O(n274), .CO(n275)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i7  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] ), 
            .I1(1'b0), .CI(n279), .O(n276), .CO(n277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i6  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] ), 
            .I1(1'b0), .CI(n281), .O(n278), .CO(n279)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i5  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] ), 
            .I1(1'b0), .CI(n283), .O(n280), .CO(n281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i4  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] ), 
            .I1(1'b0), .CI(n285), .O(n282), .CO(n283)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i3  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] ), 
            .I1(1'b0), .CI(n759), .O(n284), .CO(n285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i9  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
            .I1(1'b0), .CI(n288), .O(n286)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i8  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] ), 
            .I1(1'b0), .CI(n290), .O(n287), .CO(n288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i7  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] ), 
            .I1(1'b0), .CI(n292), .O(n289), .CO(n290)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i6  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] ), 
            .I1(1'b0), .CI(n294), .O(n291), .CO(n292)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i5  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] ), 
            .I1(1'b0), .CI(n296), .O(n293), .CO(n294)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i4  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] ), 
            .I1(1'b0), .CI(n755), .O(n295), .CO(n296)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i9  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11] ), 
            .I1(n1553), .CI(n299), .O(n297)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i8  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10] ), 
            .I1(n1556), .CI(n301), .O(n298), .CO(n299)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i7  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9] ), 
            .I1(n1559), .CI(n303), .O(n300), .CO(n301)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i6  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] ), 
            .I1(n1562), .CI(n305), .CO(n303)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i5  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] ), 
            .I1(n1565), .CI(n307), .CO(n305)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i4  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] ), 
            .I1(n1568), .CI(n309), .CO(n307)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i3  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] ), 
            .I1(n1571), .CI(n311), .CO(n309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i2  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] ), 
            .I1(n1574), .CI(n613), .CO(n311)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i14  (.I0(1'b0), 
            .I1(1'b1), .CI(n314), .O(n312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i13  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[12] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[9] ), 
            .CI(n316), .O(n313), .CO(n314)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i13 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i12  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[11] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] ), .CI(n318), 
            .O(n315), .CO(n316)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i12 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i11  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[10] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] ), .CI(n320), 
            .O(n317), .CO(n318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i11 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i10  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[9] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] ), .CI(n322), 
            .O(n319), .CO(n320)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i10 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i9  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] ), .CI(n324), 
            .O(n321), .CO(n322)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i8  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] ), .CI(n326), 
            .O(n323), .CO(n324)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i7  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] ), .CI(n328), 
            .O(n325), .CO(n326)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i6  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] ), .CI(n330), 
            .O(n327), .CO(n328)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] ), .CI(n602), 
            .O(n329), .CO(n330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i10  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[9] ), 
            .I1(1'b0), .CI(n333), .O(n331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i10 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i9  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] ), 
            .I1(1'b0), .CI(n335), .O(n332), .CO(n333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i8  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] ), 
            .I1(1'b0), .CI(n337), .O(n334), .CO(n335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i7  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] ), 
            .I1(1'b0), .CI(n339), .O(n336), .CO(n337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i6  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] ), 
            .I1(1'b0), .CI(n341), .O(n338), .CO(n339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i5  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] ), 
            .I1(1'b0), .CI(n343), .O(n340), .CO(n341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i4  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] ), 
            .I1(1'b0), .CI(n345), .O(n342), .CO(n343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i3  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] ), 
            .I1(1'b0), .CI(n598), .O(n344), .CO(n345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i13  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12] ), 
            .I1(1'b0), .CI(n382), .O(n380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i13 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i12  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] ), 
            .I1(1'b0), .CI(n398), .O(n381), .CO(n382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i12 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i11  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] ), 
            .I1(1'b0), .CI(n406), .O(n397), .CO(n398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i11 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/sub_21/add_2/i2  (.I0(\u_axi4_ctrl/wfifo_cnt[1] ), 
            .I1(1'b1), .CI(n517), .O(n399), .CO(n400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(90)
    defparam \u_axi4_ctrl/sub_21/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/sub_21/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i2  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] ), .CI(1'b0), 
            .O(n401), .CO(n402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i10  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] ), 
            .I1(1'b0), .CI(n410), .O(n405), .CO(n406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i10 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i9  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] ), 
            .I1(1'b0), .CI(n414), .O(n409), .CO(n410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_104/i2  (.I0(\u_axi4_ctrl/awaddr[11] ), .I1(\u_axi4_ctrl/awaddr[10] ), 
            .CI(1'b0), .O(n411), .CO(n412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(294)
    defparam \u_axi4_ctrl/add_104/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_104/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i8  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] ), 
            .I1(1'b0), .CI(n416), .O(n413), .CO(n414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i7  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] ), 
            .I1(1'b0), .CI(n419), .O(n415), .CO(n416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i6  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] ), 
            .I1(1'b0), .CI(n421), .O(n418), .CO(n419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i5  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] ), 
            .I1(1'b0), .CI(n423), .O(n420), .CO(n421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i4  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] ), 
            .I1(1'b0), .CI(n570), .O(n422), .CO(n423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_130/i14  (.I0(\u_axi4_ctrl/araddr[23] ), .I1(1'b0), 
            .CI(n427), .O(n425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(311)
    defparam \u_axi4_ctrl/add_130/i14 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_130/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_130/i13  (.I0(\u_axi4_ctrl/araddr[22] ), .I1(1'b0), 
            .CI(n481), .O(n426), .CO(n427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(311)
    defparam \u_axi4_ctrl/add_130/i13 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_130/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_130/i2  (.I0(\u_axi4_ctrl/araddr[11] ), .I1(\u_axi4_ctrl/araddr[10] ), 
            .CI(1'b0), .O(n460), .CO(n461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(311)
    defparam \u_axi4_ctrl/add_130/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_130/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_130/i3  (.I0(\u_axi4_ctrl/araddr[12] ), .I1(1'b0), 
            .CI(n461), .O(n470), .CO(n471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(311)
    defparam \u_axi4_ctrl/add_130/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_130/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_130/i12  (.I0(\u_axi4_ctrl/araddr[21] ), .I1(1'b0), 
            .CI(n483), .O(n480), .CO(n481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(311)
    defparam \u_axi4_ctrl/add_130/i12 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_130/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_130/i11  (.I0(\u_axi4_ctrl/araddr[20] ), .I1(1'b0), 
            .CI(n485), .O(n482), .CO(n483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(311)
    defparam \u_axi4_ctrl/add_130/i11 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_130/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_130/i10  (.I0(\u_axi4_ctrl/araddr[19] ), .I1(1'b0), 
            .CI(n487), .O(n484), .CO(n485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(311)
    defparam \u_axi4_ctrl/add_130/i10 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_130/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_130/i9  (.I0(\u_axi4_ctrl/araddr[18] ), .I1(1'b0), 
            .CI(n489), .O(n486), .CO(n487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(311)
    defparam \u_axi4_ctrl/add_130/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_130/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_130/i8  (.I0(\u_axi4_ctrl/araddr[17] ), .I1(1'b0), 
            .CI(n491), .O(n488), .CO(n489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(311)
    defparam \u_axi4_ctrl/add_130/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_130/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_130/i7  (.I0(\u_axi4_ctrl/araddr[16] ), .I1(1'b0), 
            .CI(n540), .O(n490), .CO(n491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(311)
    defparam \u_axi4_ctrl/add_130/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_130/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/sub_21/add_2/i1  (.I0(\u_axi4_ctrl/wfifo_cnt[0] ), 
            .I1(1'b0), .CI(n2553), .O(n516), .CO(n517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(90)
    defparam \u_axi4_ctrl/sub_21/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/sub_21/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_130/i6  (.I0(\u_axi4_ctrl/araddr[15] ), .I1(1'b0), 
            .CI(n542), .O(n539), .CO(n540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(311)
    defparam \u_axi4_ctrl/add_130/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_130/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_130/i5  (.I0(\u_axi4_ctrl/araddr[14] ), .I1(1'b0), 
            .CI(n544), .O(n541), .CO(n542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(311)
    defparam \u_axi4_ctrl/add_130/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_130/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_130/i4  (.I0(\u_axi4_ctrl/araddr[13] ), .I1(1'b0), 
            .CI(n471), .O(n543), .CO(n544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(311)
    defparam \u_axi4_ctrl/add_130/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_130/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_104/i14  (.I0(\u_axi4_ctrl/awaddr[23] ), .I1(1'b0), 
            .CI(n553), .O(n551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(294)
    defparam \u_axi4_ctrl/add_104/i14 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_104/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_104/i13  (.I0(\u_axi4_ctrl/awaddr[22] ), .I1(1'b0), 
            .CI(n555), .O(n552), .CO(n553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(294)
    defparam \u_axi4_ctrl/add_104/i13 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_104/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_104/i12  (.I0(\u_axi4_ctrl/awaddr[21] ), .I1(1'b0), 
            .CI(n560), .O(n554), .CO(n555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(294)
    defparam \u_axi4_ctrl/add_104/i12 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_104/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_104/i11  (.I0(\u_axi4_ctrl/awaddr[20] ), .I1(1'b0), 
            .CI(n564), .O(n559), .CO(n560)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(294)
    defparam \u_axi4_ctrl/add_104/i11 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_104/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_104/i10  (.I0(\u_axi4_ctrl/awaddr[19] ), .I1(1'b0), 
            .CI(n566), .O(n563), .CO(n564)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(294)
    defparam \u_axi4_ctrl/add_104/i10 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_104/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_104/i9  (.I0(\u_axi4_ctrl/awaddr[18] ), .I1(1'b0), 
            .CI(n594), .O(n565), .CO(n566)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(294)
    defparam \u_axi4_ctrl/add_104/i9 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_104/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i3  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] ), 
            .I1(1'b0), .CI(n402), .O(n569), .CO(n570)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_42/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_104/i8  (.I0(\u_axi4_ctrl/awaddr[17] ), .I1(1'b0), 
            .CI(n714), .O(n593), .CO(n594)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(294)
    defparam \u_axi4_ctrl/add_104/i8 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_104/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i2  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] ), .CI(1'b0), 
            .O(n597), .CO(n598)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_46/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i4  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] ), .CI(n2554), 
            .O(n601), .CO(n602)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i1  (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] ), 
            .I1(n1776), .CI(n2555), .CO(n613)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_104/i7  (.I0(\u_axi4_ctrl/awaddr[16] ), .I1(1'b0), 
            .CI(n716), .O(n713), .CO(n714)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(294)
    defparam \u_axi4_ctrl/add_104/i7 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_104/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_104/i6  (.I0(\u_axi4_ctrl/awaddr[15] ), .I1(1'b0), 
            .CI(n718), .O(n715), .CO(n716)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(294)
    defparam \u_axi4_ctrl/add_104/i6 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_104/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_104/i5  (.I0(\u_axi4_ctrl/awaddr[14] ), .I1(1'b0), 
            .CI(n720), .O(n717), .CO(n718)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(294)
    defparam \u_axi4_ctrl/add_104/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_104/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_104/i4  (.I0(\u_axi4_ctrl/awaddr[13] ), .I1(1'b0), 
            .CI(n722), .O(n719), .CO(n720)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(294)
    defparam \u_axi4_ctrl/add_104/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_104/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/add_104/i3  (.I0(\u_axi4_ctrl/awaddr[12] ), .I1(1'b0), 
            .CI(n412), .O(n721), .CO(n722)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(294)
    defparam \u_axi4_ctrl/add_104/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/add_104/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/sub_21/add_2/i5  (.I0(\u_axi4_ctrl/wfifo_cnt[4] ), 
            .I1(1'b1), .CI(n725), .O(n723)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(90)
    defparam \u_axi4_ctrl/sub_21/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/sub_21/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/sub_21/add_2/i4  (.I0(\u_axi4_ctrl/wfifo_cnt[3] ), 
            .I1(1'b1), .CI(n727), .O(n724), .CO(n725)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(90)
    defparam \u_axi4_ctrl/sub_21/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/sub_21/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/sub_21/add_2/i3  (.I0(\u_axi4_ctrl/wfifo_cnt[2] ), 
            .I1(1'b1), .CI(n400), .O(n726), .CO(n727)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(90)
    defparam \u_axi4_ctrl/sub_21/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/sub_21/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_39/i10  (.I0(\u_VsyHsyGenerator/frameCnt_value[9] ), 
            .I1(1'b0), .CI(n767), .O(n728)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(158)
    defparam \u_VsyHsyGenerator/add_39/i10 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_39/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i2  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] ), .CI(1'b0), 
            .O(n747), .CO(n748)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i3  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] ), 
            .I1(1'b0), .CI(n748), .O(n754), .CO(n755)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1272)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i3 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_44/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i2  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] ), .CI(1'b0), 
            .O(n758), .CO(n759)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1282)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i2 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/add_48/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i1  (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] ), 
            .CI(n2556), .O(n761), .CO(n762)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \u_VsyHsyGenerator/add_39/i9  (.I0(\u_VsyHsyGenerator/frameCnt_value[8] ), 
            .I1(1'b0), .CI(n870), .O(n766), .CO(n767)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(158)
    defparam \u_VsyHsyGenerator/add_39/i9 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_39/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_7/i2  (.I0(\u_lcd_driver/hcnt[1] ), .I1(\u_lcd_driver/hcnt[0] ), 
            .CI(1'b0), .O(n776), .CO(n777)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(72)
    defparam \u_lcd_driver/add_7/i2 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_7/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_39/i8  (.I0(\u_VsyHsyGenerator/frameCnt_value[7] ), 
            .I1(1'b0), .CI(n889), .O(n869), .CO(n870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(158)
    defparam \u_VsyHsyGenerator/add_39/i8 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_39/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_39/i7  (.I0(\u_VsyHsyGenerator/frameCnt_value[6] ), 
            .I1(1'b0), .CI(n891), .O(n888), .CO(n889)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(158)
    defparam \u_VsyHsyGenerator/add_39/i7 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_39/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_39/i6  (.I0(\u_VsyHsyGenerator/frameCnt_value[5] ), 
            .I1(1'b0), .CI(n893), .O(n890), .CO(n891)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(158)
    defparam \u_VsyHsyGenerator/add_39/i6 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_39/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_39/i5  (.I0(\u_VsyHsyGenerator/frameCnt_value[4] ), 
            .I1(1'b0), .CI(n895), .O(n892), .CO(n893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(158)
    defparam \u_VsyHsyGenerator/add_39/i5 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_39/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_39/i4  (.I0(\u_VsyHsyGenerator/frameCnt_value[3] ), 
            .I1(1'b0), .CI(n897), .O(n894), .CO(n895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(158)
    defparam \u_VsyHsyGenerator/add_39/i4 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_39/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_39/i3  (.I0(\u_VsyHsyGenerator/frameCnt_value[2] ), 
            .I1(1'b0), .CI(n899), .O(n896), .CO(n897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(158)
    defparam \u_VsyHsyGenerator/add_39/i3 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_39/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_39/i2  (.I0(\u_VsyHsyGenerator/frameCnt_value[1] ), 
            .I1(1'b0), .CI(n201), .O(n898), .CO(n899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(158)
    defparam \u_VsyHsyGenerator/add_39/i2 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_39/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_31/i11  (.I0(\u_VsyHsyGenerator/pCnt_value[10] ), 
            .I1(1'b0), .CI(n902), .O(n900)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(129)
    defparam \u_VsyHsyGenerator/add_31/i11 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_31/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_31/i10  (.I0(\u_VsyHsyGenerator/pCnt_value[9] ), 
            .I1(1'b0), .CI(n904), .O(n901), .CO(n902)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(129)
    defparam \u_VsyHsyGenerator/add_31/i10 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_31/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_31/i9  (.I0(\u_VsyHsyGenerator/pCnt_value[8] ), 
            .I1(1'b0), .CI(n906), .O(n903), .CO(n904)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(129)
    defparam \u_VsyHsyGenerator/add_31/i9 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_31/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_31/i8  (.I0(\u_VsyHsyGenerator/pCnt_value[7] ), 
            .I1(1'b0), .CI(n908), .O(n905), .CO(n906)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(129)
    defparam \u_VsyHsyGenerator/add_31/i8 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_31/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_31/i7  (.I0(\u_VsyHsyGenerator/pCnt_value[6] ), 
            .I1(1'b0), .CI(n910), .O(n907), .CO(n908)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(129)
    defparam \u_VsyHsyGenerator/add_31/i7 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_31/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_31/i6  (.I0(\u_VsyHsyGenerator/pCnt_value[5] ), 
            .I1(1'b0), .CI(n912), .O(n909), .CO(n910)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(129)
    defparam \u_VsyHsyGenerator/add_31/i6 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_31/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_31/i5  (.I0(\u_VsyHsyGenerator/pCnt_value[4] ), 
            .I1(1'b0), .CI(n914), .O(n911), .CO(n912)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(129)
    defparam \u_VsyHsyGenerator/add_31/i5 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_31/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_31/i4  (.I0(\u_VsyHsyGenerator/pCnt_value[3] ), 
            .I1(1'b0), .CI(n916), .O(n913), .CO(n914)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(129)
    defparam \u_VsyHsyGenerator/add_31/i4 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_31/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_31/i3  (.I0(\u_VsyHsyGenerator/pCnt_value[2] ), 
            .I1(1'b0), .CI(n918), .O(n915), .CO(n916)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(129)
    defparam \u_VsyHsyGenerator/add_31/i3 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_31/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_31/i2  (.I0(\u_VsyHsyGenerator/pCnt_value[1] ), 
            .I1(1'b0), .CI(n199), .O(n917), .CO(n918)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(129)
    defparam \u_VsyHsyGenerator/add_31/i2 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_31/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_24/i10  (.I0(\u_VsyHsyGenerator/hsynCnt_value[9] ), 
            .I1(1'b0), .CI(n921), .O(n919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(102)
    defparam \u_VsyHsyGenerator/add_24/i10 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_24/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_24/i9  (.I0(\u_VsyHsyGenerator/hsynCnt_value[8] ), 
            .I1(1'b0), .CI(n923), .O(n920), .CO(n921)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(102)
    defparam \u_VsyHsyGenerator/add_24/i9 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_24/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_24/i8  (.I0(\u_VsyHsyGenerator/hsynCnt_value[7] ), 
            .I1(1'b0), .CI(n925), .O(n922), .CO(n923)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(102)
    defparam \u_VsyHsyGenerator/add_24/i8 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_24/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_24/i7  (.I0(\u_VsyHsyGenerator/hsynCnt_value[6] ), 
            .I1(1'b0), .CI(n927), .O(n924), .CO(n925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(102)
    defparam \u_VsyHsyGenerator/add_24/i7 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_24/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_24/i6  (.I0(\u_VsyHsyGenerator/hsynCnt_value[5] ), 
            .I1(1'b0), .CI(n929), .O(n926), .CO(n927)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(102)
    defparam \u_VsyHsyGenerator/add_24/i6 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_24/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_24/i5  (.I0(\u_VsyHsyGenerator/hsynCnt_value[4] ), 
            .I1(1'b0), .CI(n931), .O(n928), .CO(n929)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(102)
    defparam \u_VsyHsyGenerator/add_24/i5 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_24/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_24/i4  (.I0(\u_VsyHsyGenerator/hsynCnt_value[3] ), 
            .I1(1'b0), .CI(n947), .O(n930), .CO(n931)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(102)
    defparam \u_VsyHsyGenerator/add_24/i4 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_24/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_24/i3  (.I0(\u_VsyHsyGenerator/hsynCnt_value[2] ), 
            .I1(1'b0), .CI(n949), .O(n946), .CO(n947)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(102)
    defparam \u_VsyHsyGenerator/add_24/i3 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_24/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \u_VsyHsyGenerator/add_24/i2  (.I0(\u_VsyHsyGenerator/hsynCnt_value[1] ), 
            .I1(1'b0), .CI(n177), .O(n948), .CO(n949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\VsyHsyGenerator.v(102)
    defparam \u_VsyHsyGenerator/add_24/i2 .I0_POLARITY = 1'b1;
    defparam \u_VsyHsyGenerator/add_24/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i20  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19] ), 
            .I1(1'b1), .CI(n952), .O(n950)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i20 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i20 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i19  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18] ), 
            .I1(1'b1), .CI(n954), .O(n951), .CO(n952)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i19 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i19 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i18  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17] ), 
            .I1(1'b1), .CI(n956), .O(n953), .CO(n954)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i18 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i18 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i17  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16] ), 
            .I1(1'b1), .CI(n958), .O(n955), .CO(n956)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i17 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i17 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i16  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15] ), 
            .I1(1'b1), .CI(n960), .O(n957), .CO(n958)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i16 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i16 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i15  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14] ), 
            .I1(1'b1), .CI(n962), .O(n959), .CO(n960)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i15 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i15 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i14  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13] ), 
            .I1(1'b1), .CI(n964), .O(n961), .CO(n962)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i14 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i14 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i13  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12] ), 
            .I1(1'b1), .CI(n966), .O(n963), .CO(n964)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i13 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i12  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11] ), 
            .I1(1'b1), .CI(n968), .O(n965), .CO(n966)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i12 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i11  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10] ), 
            .I1(1'b1), .CI(n970), .O(n967), .CO(n968)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i10  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9] ), 
            .I1(1'b1), .CI(n972), .O(n969), .CO(n970)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i9  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8] ), 
            .I1(1'b1), .CI(n990), .O(n971), .CO(n972)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i8  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7] ), 
            .I1(1'b1), .CI(n1007), .O(n989), .CO(n990)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i7  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6] ), 
            .I1(1'b1), .CI(n1009), .O(n1006), .CO(n1007)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i6  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5] ), 
            .I1(1'b1), .CI(n1141), .O(n1008), .CO(n1009)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \u_lcd_driver/add_17/i2  (.I0(\u_lcd_driver/vcnt[1] ), .I1(\u_lcd_driver/vcnt[0] ), 
            .CI(1'b0), .O(n1137), .CO(n1138)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\lcd_driver.v(89)
    defparam \u_lcd_driver/add_17/i2 .I0_POLARITY = 1'b1;
    defparam \u_lcd_driver/add_17/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i5  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4] ), 
            .I1(1'b1), .CI(n1143), .O(n1140), .CO(n1141)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i4  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3] ), 
            .I1(1'b1), .CI(n1157), .O(n1142), .CO(n1143)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i3  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2] ), 
            .I1(1'b1), .CI(n1159), .O(n1156), .CO(n1157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i2  (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1] ), 
            .I1(1'b1), .CI(n163), .O(n1158), .CO(n1159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \add_7/i8  (.I0(\PowerOnResetCnt[7] ), .I1(1'b0), .CI(n1162), 
            .O(n1160)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(98)
    defparam \add_7/i8 .I0_POLARITY = 1'b1;
    defparam \add_7/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \add_7/i7  (.I0(\PowerOnResetCnt[6] ), .I1(1'b0), .CI(n1164), 
            .O(n1161), .CO(n1162)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(98)
    defparam \add_7/i7 .I0_POLARITY = 1'b1;
    defparam \add_7/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \add_7/i6  (.I0(\PowerOnResetCnt[5] ), .I1(1'b0), .CI(n1166), 
            .O(n1163), .CO(n1164)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(98)
    defparam \add_7/i6 .I0_POLARITY = 1'b1;
    defparam \add_7/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \add_7/i5  (.I0(\PowerOnResetCnt[4] ), .I1(1'b0), .CI(n1168), 
            .O(n1165), .CO(n1166)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(98)
    defparam \add_7/i5 .I0_POLARITY = 1'b1;
    defparam \add_7/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \add_7/i4  (.I0(\PowerOnResetCnt[3] ), .I1(1'b0), .CI(n1170), 
            .O(n1167), .CO(n1168)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(98)
    defparam \add_7/i4 .I0_POLARITY = 1'b1;
    defparam \add_7/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \add_7/i3  (.I0(\PowerOnResetCnt[2] ), .I1(1'b0), .CI(n1172), 
            .O(n1169), .CO(n1170)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(98)
    defparam \add_7/i3 .I0_POLARITY = 1'b1;
    defparam \add_7/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \add_7/i2  (.I0(\PowerOnResetCnt[1] ), .I1(1'b0), .CI(n1174), 
            .O(n1171), .CO(n1172)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(98)
    defparam \add_7/i2 .I0_POLARITY = 1'b1;
    defparam \add_7/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \add_7/i1  (.I0(\PowerOnResetCnt[0] ), .I1(\reduce_nand_6/n7 ), 
            .CI(1'b0), .O(n1173), .CO(n1174)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\T35_Sensor_DDR3_LCD_Test.v(98)
    defparam \add_7/i1 .I0_POLARITY = 1'b1;
    defparam \add_7/i1 .I1_POLARITY = 1'b0;
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12  (.WCLK(\clk_12M_i~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\XYCrop_frame_Gray[15] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[7], 
            DdrCtrl_WDATA_0[23], DdrCtrl_WDATA_0[39], DdrCtrl_WDATA_0[55], 
            DdrCtrl_WDATA_0[71], DdrCtrl_WDATA_0[87], DdrCtrl_WDATA_0[103], 
            DdrCtrl_WDATA_0[119]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=8, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .READ_WIDTH = 8;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12  (.WCLK(\clk_12M_i~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\XYCrop_frame_Gray[14] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[13], 
            DdrCtrl_WDATA_0[29], DdrCtrl_WDATA_0[45], DdrCtrl_WDATA_0[61], 
            DdrCtrl_WDATA_0[77], DdrCtrl_WDATA_0[93], DdrCtrl_WDATA_0[109], 
            DdrCtrl_WDATA_0[125]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=8, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .READ_WIDTH = 8;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$m12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12  (.WCLK(\clk_12M_i~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\XYCrop_frame_Gray[15] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[12], 
            DdrCtrl_WDATA_0[28], DdrCtrl_WDATA_0[44], DdrCtrl_WDATA_0[60], 
            DdrCtrl_WDATA_0[76], DdrCtrl_WDATA_0[92], DdrCtrl_WDATA_0[108], 
            DdrCtrl_WDATA_0[124]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=8, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .READ_WIDTH = 8;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$l12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12  (.WCLK(\clk_12M_i~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\XYCrop_frame_Gray[14] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[11], 
            DdrCtrl_WDATA_0[27], DdrCtrl_WDATA_0[43], DdrCtrl_WDATA_0[59], 
            DdrCtrl_WDATA_0[75], DdrCtrl_WDATA_0[91], DdrCtrl_WDATA_0[107], 
            DdrCtrl_WDATA_0[123]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=8, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .READ_WIDTH = 8;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$k12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1  (.WCLK(\clk_12M_i~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\XYCrop_frame_Gray[15] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[15], 
            DdrCtrl_WDATA_0[31], DdrCtrl_WDATA_0[47], DdrCtrl_WDATA_0[63], 
            DdrCtrl_WDATA_0[79], DdrCtrl_WDATA_0[95], DdrCtrl_WDATA_0[111], 
            DdrCtrl_WDATA_0[127]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=8, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .READ_WIDTH = 8;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$o1 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2  (.WCLK(\clk_12M_i~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\XYCrop_frame_Gray[9] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[0], 
            DdrCtrl_WDATA_0[16], DdrCtrl_WDATA_0[32], DdrCtrl_WDATA_0[48], 
            DdrCtrl_WDATA_0[64], DdrCtrl_WDATA_0[80], DdrCtrl_WDATA_0[96], 
            DdrCtrl_WDATA_0[112]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=8, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .READ_WIDTH = 8;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12  (.WCLK(\clk_12M_i~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\XYCrop_frame_Gray[9] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[6], 
            DdrCtrl_WDATA_0[22], DdrCtrl_WDATA_0[38], DdrCtrl_WDATA_0[54], 
            DdrCtrl_WDATA_0[70], DdrCtrl_WDATA_0[86], DdrCtrl_WDATA_0[102], 
            DdrCtrl_WDATA_0[118]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=8, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .READ_WIDTH = 8;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12  (.WCLK(\clk_12M_i~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\XYCrop_frame_Gray[15] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[10], 
            DdrCtrl_WDATA_0[26], DdrCtrl_WDATA_0[42], DdrCtrl_WDATA_0[58], 
            DdrCtrl_WDATA_0[74], DdrCtrl_WDATA_0[90], DdrCtrl_WDATA_0[106], 
            DdrCtrl_WDATA_0[122]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=8, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .READ_WIDTH = 8;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$j12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12  (.WCLK(\clk_12M_i~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\XYCrop_frame_Gray[5] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[5], 
            DdrCtrl_WDATA_0[21], DdrCtrl_WDATA_0[37], DdrCtrl_WDATA_0[53], 
            DdrCtrl_WDATA_0[69], DdrCtrl_WDATA_0[85], DdrCtrl_WDATA_0[101], 
            DdrCtrl_WDATA_0[117]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=8, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .READ_WIDTH = 8;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12  (.WCLK(\clk_12M_i~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\XYCrop_frame_Gray[9] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[9], 
            DdrCtrl_WDATA_0[25], DdrCtrl_WDATA_0[41], DdrCtrl_WDATA_0[57], 
            DdrCtrl_WDATA_0[73], DdrCtrl_WDATA_0[89], DdrCtrl_WDATA_0[105], 
            DdrCtrl_WDATA_0[121]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=8, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .READ_WIDTH = 8;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$i12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12  (.WCLK(\clk_12M_i~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\XYCrop_frame_Gray[5] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[4], 
            DdrCtrl_WDATA_0[20], DdrCtrl_WDATA_0[36], DdrCtrl_WDATA_0[52], 
            DdrCtrl_WDATA_0[68], DdrCtrl_WDATA_0[84], DdrCtrl_WDATA_0[100], 
            DdrCtrl_WDATA_0[116]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=8, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .READ_WIDTH = 8;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12  (.WCLK(\clk_12M_i~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\XYCrop_frame_Gray[14] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[3], 
            DdrCtrl_WDATA_0[19], DdrCtrl_WDATA_0[35], DdrCtrl_WDATA_0[51], 
            DdrCtrl_WDATA_0[67], DdrCtrl_WDATA_0[83], DdrCtrl_WDATA_0[99], 
            DdrCtrl_WDATA_0[115]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=8, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .READ_WIDTH = 8;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12  (.WCLK(\clk_12M_i~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\XYCrop_frame_Gray[14] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[14], 
            DdrCtrl_WDATA_0[30], DdrCtrl_WDATA_0[46], DdrCtrl_WDATA_0[62], 
            DdrCtrl_WDATA_0[78], DdrCtrl_WDATA_0[94], DdrCtrl_WDATA_0[110], 
            DdrCtrl_WDATA_0[126]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=8, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .READ_WIDTH = 8;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$n12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\tx_slowclk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[1] , 
            \u_axi4_ctrl/rfifo_wdata[0] , \u_axi4_ctrl/rfifo_wdata[17] , 
            \u_axi4_ctrl/rfifo_wdata[16] , \u_axi4_ctrl/rfifo_wdata[33] , 
            \u_axi4_ctrl/rfifo_wdata[32] , \u_axi4_ctrl/rfifo_wdata[49] , 
            \u_axi4_ctrl/rfifo_wdata[48] , \u_axi4_ctrl/rfifo_wdata[65] , 
            \u_axi4_ctrl/rfifo_wdata[64] , \u_axi4_ctrl/rfifo_wdata[81] , 
            \u_axi4_ctrl/rfifo_wdata[80] , \u_axi4_ctrl/rfifo_wdata[97] , 
            \u_axi4_ctrl/rfifo_wdata[96] , \u_axi4_ctrl/rfifo_wdata[113] , 
            \u_axi4_ctrl/rfifo_wdata[112] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({\lcd_data[1] , \lcd_data[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .READ_WIDTH = 2;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$2 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12  (.WCLK(\clk_12M_i~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\XYCrop_frame_Gray[14] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[2], 
            DdrCtrl_WDATA_0[18], DdrCtrl_WDATA_0[34], DdrCtrl_WDATA_0[50], 
            DdrCtrl_WDATA_0[66], DdrCtrl_WDATA_0[82], DdrCtrl_WDATA_0[98], 
            DdrCtrl_WDATA_0[114]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=8, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .READ_WIDTH = 8;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12  (.WCLK(\clk_12M_i~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\XYCrop_frame_Gray[5] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[1], 
            DdrCtrl_WDATA_0[17], DdrCtrl_WDATA_0[33], DdrCtrl_WDATA_0[49], 
            DdrCtrl_WDATA_0[65], DdrCtrl_WDATA_0[81], DdrCtrl_WDATA_0[97], 
            DdrCtrl_WDATA_0[113]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=8, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .READ_WIDTH = 8;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\tx_slowclk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[5] , 
            \u_axi4_ctrl/rfifo_wdata[4] , \u_axi4_ctrl/rfifo_wdata[21] , 
            \u_axi4_ctrl/rfifo_wdata[20] , \u_axi4_ctrl/rfifo_wdata[37] , 
            \u_axi4_ctrl/rfifo_wdata[36] , \u_axi4_ctrl/rfifo_wdata[53] , 
            \u_axi4_ctrl/rfifo_wdata[52] , \u_axi4_ctrl/rfifo_wdata[69] , 
            \u_axi4_ctrl/rfifo_wdata[68] , \u_axi4_ctrl/rfifo_wdata[85] , 
            \u_axi4_ctrl/rfifo_wdata[84] , \u_axi4_ctrl/rfifo_wdata[101] , 
            \u_axi4_ctrl/rfifo_wdata[100] , \u_axi4_ctrl/rfifo_wdata[117] , 
            \u_axi4_ctrl/rfifo_wdata[116] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({\lcd_data[5] , \lcd_data[4] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .READ_WIDTH = 2;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$b12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12  (.WCLK(\clk_12M_i~O ), 
            .RCLK(\Axi_Clk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\XYCrop_frame_Gray[14] }), 
            .WADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[2] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[1] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[0] }), 
            .RADDR({\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] , \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] , 
            \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] }), .RDATA({DdrCtrl_WDATA_0[8], 
            DdrCtrl_WDATA_0[24], DdrCtrl_WDATA_0[40], DdrCtrl_WDATA_0[56], 
            DdrCtrl_WDATA_0[72], DdrCtrl_WDATA_0[88], DdrCtrl_WDATA_0[104], 
            DdrCtrl_WDATA_0[120]})) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=8, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .READ_WIDTH = 8;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .WRITE_WIDTH = 1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$h12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\tx_slowclk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[7] , 
            \u_axi4_ctrl/rfifo_wdata[6] , \u_axi4_ctrl/rfifo_wdata[23] , 
            \u_axi4_ctrl/rfifo_wdata[22] , \u_axi4_ctrl/rfifo_wdata[39] , 
            \u_axi4_ctrl/rfifo_wdata[38] , \u_axi4_ctrl/rfifo_wdata[55] , 
            \u_axi4_ctrl/rfifo_wdata[54] , \u_axi4_ctrl/rfifo_wdata[71] , 
            \u_axi4_ctrl/rfifo_wdata[70] , \u_axi4_ctrl/rfifo_wdata[87] , 
            \u_axi4_ctrl/rfifo_wdata[86] , \u_axi4_ctrl/rfifo_wdata[103] , 
            \u_axi4_ctrl/rfifo_wdata[102] , \u_axi4_ctrl/rfifo_wdata[119] , 
            \u_axi4_ctrl/rfifo_wdata[118] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({\lcd_data[7] , \lcd_data[6] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .READ_WIDTH = 2;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$c12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\tx_slowclk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[11] , 
            \u_axi4_ctrl/rfifo_wdata[10] , \u_axi4_ctrl/rfifo_wdata[27] , 
            \u_axi4_ctrl/rfifo_wdata[26] , \u_axi4_ctrl/rfifo_wdata[43] , 
            \u_axi4_ctrl/rfifo_wdata[42] , \u_axi4_ctrl/rfifo_wdata[59] , 
            \u_axi4_ctrl/rfifo_wdata[58] , \u_axi4_ctrl/rfifo_wdata[75] , 
            \u_axi4_ctrl/rfifo_wdata[74] , \u_axi4_ctrl/rfifo_wdata[91] , 
            \u_axi4_ctrl/rfifo_wdata[90] , \u_axi4_ctrl/rfifo_wdata[107] , 
            \u_axi4_ctrl/rfifo_wdata[106] , \u_axi4_ctrl/rfifo_wdata[123] , 
            \u_axi4_ctrl/rfifo_wdata[122] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({\lcd_data[11] , \lcd_data[10] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .READ_WIDTH = 2;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$e12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\tx_slowclk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[13] , 
            \u_axi4_ctrl/rfifo_wdata[12] , \u_axi4_ctrl/rfifo_wdata[29] , 
            \u_axi4_ctrl/rfifo_wdata[28] , \u_axi4_ctrl/rfifo_wdata[45] , 
            \u_axi4_ctrl/rfifo_wdata[44] , \u_axi4_ctrl/rfifo_wdata[61] , 
            \u_axi4_ctrl/rfifo_wdata[60] , \u_axi4_ctrl/rfifo_wdata[77] , 
            \u_axi4_ctrl/rfifo_wdata[76] , \u_axi4_ctrl/rfifo_wdata[93] , 
            \u_axi4_ctrl/rfifo_wdata[92] , \u_axi4_ctrl/rfifo_wdata[109] , 
            \u_axi4_ctrl/rfifo_wdata[108] , \u_axi4_ctrl/rfifo_wdata[125] , 
            \u_axi4_ctrl/rfifo_wdata[124] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({\lcd_data[13] , \lcd_data[12] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .READ_WIDTH = 2;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$f12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\tx_slowclk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[15] , 
            \u_axi4_ctrl/rfifo_wdata[14] , \u_axi4_ctrl/rfifo_wdata[31] , 
            \u_axi4_ctrl/rfifo_wdata[30] , \u_axi4_ctrl/rfifo_wdata[47] , 
            \u_axi4_ctrl/rfifo_wdata[46] , \u_axi4_ctrl/rfifo_wdata[63] , 
            \u_axi4_ctrl/rfifo_wdata[62] , \u_axi4_ctrl/rfifo_wdata[79] , 
            \u_axi4_ctrl/rfifo_wdata[78] , \u_axi4_ctrl/rfifo_wdata[95] , 
            \u_axi4_ctrl/rfifo_wdata[94] , \u_axi4_ctrl/rfifo_wdata[111] , 
            \u_axi4_ctrl/rfifo_wdata[110] , \u_axi4_ctrl/rfifo_wdata[127] , 
            \u_axi4_ctrl/rfifo_wdata[126] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({\lcd_data[15] , \lcd_data[14] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .READ_WIDTH = 2;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$g1 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\tx_slowclk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[9] , 
            \u_axi4_ctrl/rfifo_wdata[8] , \u_axi4_ctrl/rfifo_wdata[25] , 
            \u_axi4_ctrl/rfifo_wdata[24] , \u_axi4_ctrl/rfifo_wdata[41] , 
            \u_axi4_ctrl/rfifo_wdata[40] , \u_axi4_ctrl/rfifo_wdata[57] , 
            \u_axi4_ctrl/rfifo_wdata[56] , \u_axi4_ctrl/rfifo_wdata[73] , 
            \u_axi4_ctrl/rfifo_wdata[72] , \u_axi4_ctrl/rfifo_wdata[89] , 
            \u_axi4_ctrl/rfifo_wdata[88] , \u_axi4_ctrl/rfifo_wdata[105] , 
            \u_axi4_ctrl/rfifo_wdata[104] , \u_axi4_ctrl/rfifo_wdata[121] , 
            \u_axi4_ctrl/rfifo_wdata[120] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({\lcd_data[9] , \lcd_data[8] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .READ_WIDTH = 2;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$d12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_RAM_5K \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12  (.WCLK(\Axi_Clk~O ), 
            .RCLK(\tx_slowclk~O ), .WCLKE(1'b1), .WE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int ), 
            .RE(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int ), .WDATA({\u_axi4_ctrl/rfifo_wdata[3] , 
            \u_axi4_ctrl/rfifo_wdata[2] , \u_axi4_ctrl/rfifo_wdata[19] , 
            \u_axi4_ctrl/rfifo_wdata[18] , \u_axi4_ctrl/rfifo_wdata[35] , 
            \u_axi4_ctrl/rfifo_wdata[34] , \u_axi4_ctrl/rfifo_wdata[51] , 
            \u_axi4_ctrl/rfifo_wdata[50] , \u_axi4_ctrl/rfifo_wdata[67] , 
            \u_axi4_ctrl/rfifo_wdata[66] , \u_axi4_ctrl/rfifo_wdata[83] , 
            \u_axi4_ctrl/rfifo_wdata[82] , \u_axi4_ctrl/rfifo_wdata[99] , 
            \u_axi4_ctrl/rfifo_wdata[98] , \u_axi4_ctrl/rfifo_wdata[115] , 
            \u_axi4_ctrl/rfifo_wdata[114] }), .WADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] }), .RADDR({\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[2] , 
            \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[1] , \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[0] }), 
            .RDATA({\lcd_data[3] , \lcd_data[2] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=16, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_UNKNOWN", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(705)
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .READ_WIDTH = 2;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WRITE_WIDTH = 16;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .OUTPUT_REG = 1'b0;
    defparam \u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ram/ram__D$12 .WRITE_MODE = "READ_UNKNOWN";
    EFX_LUT4 LUT__3687 (.I0(\u_axi4_ctrl/state[0] ), .I1(DdrCtrl_BREADY_0), 
            .O(DdrCtrl_WVALID_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3687.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3688 (.I0(\u_axi4_ctrl/wdata_cnt_dly[0] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[1] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[2] ), .I3(\u_axi4_ctrl/wdata_cnt_dly[3] ), 
            .O(n2429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3688.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3689 (.I0(\u_axi4_ctrl/wdata_cnt_dly[0] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[1] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[2] ), .I3(\u_axi4_ctrl/wdata_cnt_dly[3] ), 
            .O(n2430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3689.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3690 (.I0(n2430), .I1(n2429), .I2(DdrCtrl_WREADY_0), 
            .O(n2431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3690.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3691 (.I0(DdrCtrl_WREADY_0), .I1(\u_axi4_ctrl/wdata_cnt_dly[4] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[5] ), .O(n2432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7e7e */ ;
    defparam LUT__3691.LUTMASK = 16'h7e7e;
    EFX_LUT4 LUT__3692 (.I0(n2432), .I1(\u_axi4_ctrl/wdata_cnt_dly[7] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[8] ), .O(n2433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__3692.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__3693 (.I0(\u_axi4_ctrl/wdata_cnt_dly[4] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[5] ), 
            .O(n2434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3693.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3694 (.I0(n2430), .I1(n2434), .I2(\u_axi4_ctrl/wdata_cnt_dly[6] ), 
            .O(\u_axi4_ctrl/n1531 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__3694.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__3695 (.I0(n2431), .I1(DdrCtrl_WVALID_0), .I2(n2433), 
            .I3(\u_axi4_ctrl/n1531 ), .O(DdrCtrl_WLAST_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__3695.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__3696 (.I0(\u_axi4_ctrl/state[1] ), .I1(\u_axi4_ctrl/state[2] ), 
            .O(n2435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3696.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3697 (.I0(n2435), .I1(\u_axi4_ctrl/state[0] ), .O(DdrCtrl_RREADY_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3697.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3698 (.I0(\u_lcd_driver/vcnt[0] ), .I1(\u_lcd_driver/vcnt[1] ), 
            .I2(\u_lcd_driver/vcnt[2] ), .O(n2436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3698.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3699 (.I0(n2436), .I1(\u_lcd_driver/vcnt[3] ), .I2(\u_lcd_driver/vcnt[4] ), 
            .I3(\u_lcd_driver/vcnt[5] ), .O(n2437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h07e0 */ ;
    defparam LUT__3699.LUTMASK = 16'h07e0;
    EFX_LUT4 LUT__3700 (.I0(\u_lcd_driver/vcnt[6] ), .I1(\u_lcd_driver/vcnt[7] ), 
            .I2(\u_lcd_driver/vcnt[8] ), .I3(\u_lcd_driver/vcnt[9] ), .O(n2438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3700.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3701 (.I0(\u_lcd_driver/vcnt[6] ), .I1(\u_lcd_driver/vcnt[9] ), 
            .I2(n2438), .I3(\u_lcd_driver/vcnt[5] ), .O(n2439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h770f */ ;
    defparam LUT__3701.LUTMASK = 16'h770f;
    EFX_LUT4 LUT__3702 (.I0(\u_lcd_driver/vcnt[7] ), .I1(\u_lcd_driver/vcnt[8] ), 
            .O(n2440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3702.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3703 (.I0(\u_lcd_driver/vcnt[10] ), .I1(\u_lcd_driver/vcnt[11] ), 
            .O(n2441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3703.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3704 (.I0(n2440), .I1(\u_lcd_driver/vcnt[9] ), .I2(\u_lcd_driver/hcnt[11] ), 
            .I3(n2441), .O(n2442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b00 */ ;
    defparam LUT__3704.LUTMASK = 16'h0b00;
    EFX_LUT4 LUT__3705 (.I0(\u_lcd_driver/hcnt[5] ), .I1(\u_lcd_driver/hcnt[6] ), 
            .I2(\u_lcd_driver/hcnt[7] ), .O(n2443)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he0e0 */ ;
    defparam LUT__3705.LUTMASK = 16'he0e0;
    EFX_LUT4 LUT__3706 (.I0(n2443), .I1(\u_lcd_driver/hcnt[8] ), .I2(\u_lcd_driver/hcnt[9] ), 
            .I3(\u_lcd_driver/hcnt[10] ), .O(n2444)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h01fe */ ;
    defparam LUT__3706.LUTMASK = 16'h01fe;
    EFX_LUT4 LUT__3707 (.I0(n2439), .I1(n2437), .I2(n2442), .I3(n2444), 
            .O(lvds_tx2_DATA[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he000 */ ;
    defparam LUT__3707.LUTMASK = 16'he000;
    EFX_LUT4 LUT__3708 (.I0(lvds_tx2_DATA[0]), .I1(\lcd_data[11] ), .O(lvds_tx0_DATA[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3708.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3709 (.I0(lvds_tx2_DATA[0]), .I1(\lcd_data[12] ), .O(lvds_tx0_DATA[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3709.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3710 (.I0(lvds_tx2_DATA[0]), .I1(\lcd_data[13] ), .O(lvds_tx0_DATA[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3710.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3711 (.I0(lvds_tx2_DATA[0]), .I1(\lcd_data[5] ), .O(lvds_tx1_DATA[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3711.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3712 (.I0(lvds_tx2_DATA[0]), .I1(\lcd_data[6] ), .O(lvds_tx1_DATA[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3712.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3713 (.I0(lvds_tx2_DATA[0]), .I1(\lcd_data[7] ), .O(lvds_tx1_DATA[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3713.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3714 (.I0(lvds_tx2_DATA[0]), .I1(\lcd_data[8] ), .O(lvds_tx1_DATA[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3714.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3715 (.I0(lvds_tx2_DATA[0]), .I1(\lcd_data[0] ), .O(lvds_tx2_DATA[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3715.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3716 (.I0(lvds_tx2_DATA[0]), .I1(\lcd_data[1] ), .O(lvds_tx2_DATA[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3716.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3717 (.I0(lvds_tx2_DATA[0]), .I1(\lcd_data[2] ), .O(lvds_tx2_DATA[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3717.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3718 (.I0(lvds_tx2_DATA[0]), .I1(\lcd_data[14] ), .O(lvds_tx3_DATA[6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3718.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3719 (.I0(lvds_tx2_DATA[0]), .I1(\lcd_data[15] ), .O(lvds_tx3_DATA[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3719.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3720 (.I0(lvds_tx2_DATA[0]), .I1(\lcd_data[9] ), .O(lvds_tx3_DATA[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3720.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3721 (.I0(lvds_tx2_DATA[0]), .I1(\lcd_data[10] ), .O(lvds_tx3_DATA[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3721.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3722 (.I0(lvds_tx2_DATA[0]), .I1(\lcd_data[3] ), .O(lvds_tx3_DATA[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3722.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3723 (.I0(lvds_tx2_DATA[0]), .I1(\lcd_data[4] ), .O(lvds_tx3_DATA[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3723.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3724 (.I0(\PowerOnResetCnt[4] ), .I1(\PowerOnResetCnt[5] ), 
            .I2(\PowerOnResetCnt[6] ), .I3(\PowerOnResetCnt[7] ), .O(n2445)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3724.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3725 (.I0(\PowerOnResetCnt[0] ), .I1(\PowerOnResetCnt[1] ), 
            .I2(\PowerOnResetCnt[2] ), .I3(\PowerOnResetCnt[3] ), .O(n2446)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3725.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3726 (.I0(n2445), .I1(n2446), .O(\reduce_nand_6/n7 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3726.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3727 (.I0(PllLocked[1]), .I1(PllLocked[0]), .O(n6_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3727.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3728 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[4] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[5] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[6] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[7] ), .O(n2447)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3728.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3729 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[0] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[1] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[2] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[3] ), .O(n2448)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3729.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3730 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[16] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[17] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[18] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[19] ), .O(n2449)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3730.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3731 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[12] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[13] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[14] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[15] ), .O(n2450)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3731.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3732 (.I0(n2447), .I1(n2448), .I2(n2449), .I3(n2450), 
            .O(n2451)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3732.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3733 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[8] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[9] ), .I2(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[10] ), 
            .I3(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt[11] ), .O(n2452)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3733.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3734 (.I0(n2451), .I1(n2452), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n15 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777 */ ;
    defparam LUT__3734.LUTMASK = 16'h7777;
    EFX_LUT4 LUT__3735 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] ), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/equal_21/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7777 */ ;
    defparam LUT__3735.LUTMASK = 16'h7777;
    EFX_LUT4 LUT__3736 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] ), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n92 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3736.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3737 (.I0(\u_VsyHsyGenerator/hsynCnt_value[3] ), .I1(\u_VsyHsyGenerator/hsynCnt_value[4] ), 
            .I2(\u_VsyHsyGenerator/hsynCnt_value[5] ), .I3(\u_VsyHsyGenerator/hsynCnt_value[6] ), 
            .O(n2453)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__3737.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__3738 (.I0(\u_VsyHsyGenerator/hsynCnt_value[7] ), .I1(\u_VsyHsyGenerator/hsynCnt_value[8] ), 
            .O(n2454)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3738.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3739 (.I0(n2454), .I1(n2453), .I2(\u_VsyHsyGenerator/hsynCnt_value[9] ), 
            .O(n2455)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__3739.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__3740 (.I0(\u_VsyHsyGenerator/vsynDl[1] ), .I1(\u_VsyHsyGenerator/vsynDl[2] ), 
            .I2(XYCrop_frame_vsync), .O(n2456)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__3740.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__3741 (.I0(\u_VsyHsyGenerator/pCnt_value[7] ), .I1(\u_VsyHsyGenerator/pCnt_value[8] ), 
            .I2(\u_VsyHsyGenerator/pCnt_value[9] ), .O(n2457)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__3741.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__3742 (.I0(\u_VsyHsyGenerator/pCnt_value[2] ), .I1(\u_VsyHsyGenerator/pCnt_value[3] ), 
            .I2(\u_VsyHsyGenerator/pCnt_value[4] ), .O(n2458)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__3742.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__3743 (.I0(\u_VsyHsyGenerator/pCntInc ), .I1(\u_VsyHsyGenerator/pCnt_value[10] ), 
            .O(n2459)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3743.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3744 (.I0(\u_VsyHsyGenerator/pCnt_value[0] ), .I1(\u_VsyHsyGenerator/pCnt_value[1] ), 
            .I2(\u_VsyHsyGenerator/pCnt_value[5] ), .I3(\u_VsyHsyGenerator/pCnt_value[6] ), 
            .O(n2460)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3744.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3745 (.I0(n2457), .I1(n2458), .I2(n2459), .I3(n2460), 
            .O(n2461)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3745.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3746 (.I0(n2455), .I1(n2456), .I2(n2461), .I3(\u_VsyHsyGenerator/vsynDl[0] ), 
            .O(\u_VsyHsyGenerator/n519 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__3746.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__3747 (.I0(\u_VsyHsyGenerator/pCnt_value[0] ), .I1(\u_VsyHsyGenerator/pCnt_value[1] ), 
            .O(n2462)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3747.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3748 (.I0(\u_VsyHsyGenerator/pCnt_value[5] ), .I1(\u_VsyHsyGenerator/pCnt_value[6] ), 
            .O(n2463)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3748.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3749 (.I0(n2462), .I1(n2457), .I2(n2463), .I3(n2458), 
            .O(n2464)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3749.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3750 (.I0(n2455), .I1(\u_VsyHsyGenerator/n519 ), .I2(n2459), 
            .I3(n2464), .O(n1405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__3750.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__3751 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[0] ), 
            .I1(\U0_DDR_Reset/u_ddr_reset_sequencer/cnt_start[1] ), .O(\U0_DDR_Reset/u_ddr_reset_sequencer/n91 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'heeee */ ;
    defparam LUT__3751.LUTMASK = 16'heeee;
    EFX_LUT4 LUT__3752 (.I0(\u_VsyHsyGenerator/hsynCnt_value[3] ), .I1(\u_VsyHsyGenerator/hsynCnt_value[4] ), 
            .I2(\u_VsyHsyGenerator/hsynCnt_value[6] ), .I3(\u_VsyHsyGenerator/hsynCnt_value[9] ), 
            .O(n2465)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3752.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3753 (.I0(\u_VsyHsyGenerator/vsynDl[0] ), .I1(\u_VsyHsyGenerator/pCnt_value[10] ), 
            .I2(n2465), .O(n2466)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3753.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3754 (.I0(\u_VsyHsyGenerator/hsynCnt_value[0] ), .I1(\u_VsyHsyGenerator/hsynCnt_value[1] ), 
            .I2(\u_VsyHsyGenerator/hsynCnt_value[2] ), .I3(\u_VsyHsyGenerator/hsynCnt_value[5] ), 
            .O(n2467)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3754.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3755 (.I0(n2454), .I1(n2467), .O(n2468)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3755.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3756 (.I0(n2466), .I1(n2464), .I2(n2455), .I3(n2468), 
            .O(n1429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf800 */ ;
    defparam LUT__3756.LUTMASK = 16'hf800;
    EFX_LUT4 LUT__3757 (.I0(\u_axi4_ctrl/state[0] ), .I1(\u_axi4_ctrl/state[2] ), 
            .I2(\u_axi4_ctrl/state[1] ), .I3(DdrCtrl_WREADY_0), .O(\u_axi4_ctrl/n370 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__3757.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__3758 (.I0(n312), .I1(n317), .I2(n321), .I3(n323), 
            .O(n2469)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3758.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3759 (.I0(n327), .I1(n329), .I2(n601), .I3(n2469), 
            .O(n2470)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3759.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3760 (.I0(n313), .I1(n315), .I2(n319), .I3(n325), 
            .O(n2471)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3760.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3761 (.I0(n2470), .I1(n2471), .O(n2472)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3761.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3762 (.I0(\u_axi4_ctrl/n370 ), .I1(\u_axi4_ctrl/wfifo_empty ), 
            .I2(n2472), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/rd_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__3762.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__3763 (.I0(\u_VsyHsyGenerator/hsynCnt_value[6] ), .I1(\u_VsyHsyGenerator/hsynCnt_value[7] ), 
            .I2(\u_VsyHsyGenerator/hsynCnt_value[8] ), .O(n2473)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__3763.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__3764 (.I0(\u_VsyHsyGenerator/hsynCnt_value[0] ), .I1(\u_VsyHsyGenerator/hsynCnt_value[2] ), 
            .I2(\u_VsyHsyGenerator/hsynCnt_value[3] ), .I3(n2473), .O(n2474)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3764.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3765 (.I0(\u_VsyHsyGenerator/hsynCnt_value[1] ), .I1(\u_VsyHsyGenerator/hsynCnt_value[2] ), 
            .I2(\u_VsyHsyGenerator/hsynCnt_value[3] ), .O(n2475)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__3765.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__3766 (.I0(n2475), .I1(\u_VsyHsyGenerator/hsynCnt_value[5] ), 
            .I2(\u_VsyHsyGenerator/hsynCnt_value[4] ), .I3(n2473), .O(n2476)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbf00 */ ;
    defparam LUT__3766.LUTMASK = 16'hbf00;
    EFX_LUT4 LUT__3767 (.I0(n2474), .I1(n2476), .I2(\u_VsyHsyGenerator/hsynCnt_value[9] ), 
            .O(n2477)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'he3e3 */ ;
    defparam LUT__3767.LUTMASK = 16'he3e3;
    EFX_LUT4 LUT__3768 (.I0(\u_VsyHsyGenerator/pCnt_value[7] ), .I1(\u_VsyHsyGenerator/pCnt_value[8] ), 
            .I2(\u_VsyHsyGenerator/pCnt_value[9] ), .O(n2478)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3768.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3769 (.I0(n2457), .I1(n2478), .I2(\u_VsyHsyGenerator/pCnt_value[5] ), 
            .I3(\u_VsyHsyGenerator/pCnt_value[6] ), .O(n2479)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5ff3 */ ;
    defparam LUT__3769.LUTMASK = 16'h5ff3;
    EFX_LUT4 LUT__3770 (.I0(\u_VsyHsyGenerator/pCnt_value[10] ), .I1(\u_VsyHsyGenerator/pCnt_value[2] ), 
            .I2(n2462), .O(n2480)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3770.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3771 (.I0(n2479), .I1(\u_VsyHsyGenerator/pCnt_value[3] ), 
            .I2(\u_VsyHsyGenerator/pCnt_value[4] ), .I3(n2480), .O(n2481)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3771.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3772 (.I0(n2463), .I1(n2458), .I2(n2478), .O(n2482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__3772.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__3773 (.I0(\u_VsyHsyGenerator/hsynCnt_value[6] ), .I1(\u_VsyHsyGenerator/hsynCnt_value[4] ), 
            .I2(\u_VsyHsyGenerator/hsynCnt_value[5] ), .I3(\u_VsyHsyGenerator/hsynCnt_value[1] ), 
            .O(n2483)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__3773.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__3774 (.I0(\u_VsyHsyGenerator/hsynCnt_value[0] ), .I1(\u_VsyHsyGenerator/hsynCnt_value[2] ), 
            .I2(\u_VsyHsyGenerator/hsynCnt_value[3] ), .I3(n2483), .O(n2484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3774.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3775 (.I0(\u_VsyHsyGenerator/pCnt_value[5] ), .I1(\u_VsyHsyGenerator/pCnt_value[6] ), 
            .O(n2485)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3775.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3776 (.I0(n2458), .I1(n2485), .I2(n2457), .I3(\u_VsyHsyGenerator/pCnt_value[10] ), 
            .O(n2486)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h004f */ ;
    defparam LUT__3776.LUTMASK = 16'h004f;
    EFX_LUT4 LUT__3777 (.I0(n2482), .I1(n2484), .I2(n2486), .O(n2487)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3777.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3778 (.I0(n2487), .I1(n2454), .I2(n2477), .I3(n2481), 
            .O(\XYCrop_frame_Gray[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf888 */ ;
    defparam LUT__3778.LUTMASK = 16'hf888;
    EFX_LUT4 LUT__3779 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[1] ), 
            .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[0] ), 
            .I3(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] ), .O(n2488)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3779.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3780 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] ), 
            .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] ), 
            .I3(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] ), .O(n2489)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3780.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3781 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] ), .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] ), 
            .I3(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9] ), 
            .O(n2490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4182 */ ;
    defparam LUT__3781.LUTMASK = 16'h4182;
    EFX_LUT4 LUT__3782 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] ), 
            .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] ), 
            .I3(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] ), .O(n2491)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3782.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3783 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[2] ), 
            .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] ), .I3(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] ), 
            .O(n2492)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3783.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3784 (.I0(n2489), .I1(n2490), .I2(n2491), .I3(n2492), 
            .O(n2493)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3784.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3785 (.I0(n2493), .I1(n2488), .I2(XYCrop_frame_href), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/wr_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__3785.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__3786 (.I0(n2461), .I1(n198), .O(\u_VsyHsyGenerator/pCnt_valueNext[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3786.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3787 (.I0(\u_VsyHsyGenerator/frameCnt_value[0] ), .I1(\u_VsyHsyGenerator/frameCnt_value[1] ), 
            .I2(\u_VsyHsyGenerator/frameCnt_value[2] ), .I3(\u_VsyHsyGenerator/frameCnt_value[3] ), 
            .O(n2494)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3787.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3788 (.I0(\u_VsyHsyGenerator/frameCnt_value[6] ), .I1(\u_VsyHsyGenerator/frameCnt_value[7] ), 
            .I2(\u_VsyHsyGenerator/frameCnt_value[8] ), .I3(\u_VsyHsyGenerator/frameCnt_value[9] ), 
            .O(n2495)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__3788.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__3789 (.I0(\u_VsyHsyGenerator/frameCnt_value[5] ), .I1(n2494), 
            .I2(\u_VsyHsyGenerator/frameCnt_value[4] ), .I3(n2495), .O(n2496)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__3789.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__3790 (.I0(n1429), .I1(n2496), .I2(n200), .O(\u_VsyHsyGenerator/frameCnt_valueNext[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__3790.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__3791 (.I0(n2496), .I1(n1429), .O(\u_VsyHsyGenerator/n402 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3791.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3792 (.I0(n1429), .I1(\u_VsyHsyGenerator/vsynDl[0] ), 
            .I2(n2456), .O(ceg_net2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3792.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3793 (.I0(\u_VsyHsyGenerator/hsynDl[0] ), .I1(\u_VsyHsyGenerator/hsynDl[2] ), 
            .I2(XYCrop_frame_href), .I3(\u_VsyHsyGenerator/hsynDl[1] ), 
            .O(\u_VsyHsyGenerator/when_MyTopLevel_l56 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4200 */ ;
    defparam LUT__3793.LUTMASK = 16'h4200;
    EFX_LUT4 LUT__3794 (.I0(n2461), .I1(\u_VsyHsyGenerator/when_MyTopLevel_l56 ), 
            .O(ceg_net5)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3794.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3795 (.I0(n1429), .I1(n176), .O(\u_VsyHsyGenerator/hsynCnt_valueNext[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3795.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3796 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[8] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] ), 
            .I2(\u_axi4_ctrl/wfifo_empty ), .O(n1553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3796.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3797 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[7] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] ), 
            .I2(\u_axi4_ctrl/wfifo_empty ), .O(n1556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3797.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3798 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[6] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] ), 
            .I2(\u_axi4_ctrl/wfifo_empty ), .O(n1559)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3798.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3799 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[5] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] ), 
            .I2(\u_axi4_ctrl/wfifo_empty ), .O(n1562)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3799.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3800 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[4] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] ), 
            .I2(\u_axi4_ctrl/wfifo_empty ), .O(n1565)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3800.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3801 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[3] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] ), 
            .I2(\u_axi4_ctrl/wfifo_empty ), .O(n1568)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3801.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3802 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[2] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[2] ), 
            .I2(\u_axi4_ctrl/wfifo_empty ), .O(n1571)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3802.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3803 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[1] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[1] ), 
            .I2(\u_axi4_ctrl/wfifo_empty ), .O(n1574)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3803.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3804 (.I0(n2461), .I1(n917), .O(\u_VsyHsyGenerator/pCnt_valueNext[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3804.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3805 (.I0(n2461), .I1(n915), .O(\u_VsyHsyGenerator/pCnt_valueNext[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3805.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3806 (.I0(n2461), .I1(n913), .O(\u_VsyHsyGenerator/pCnt_valueNext[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3806.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3807 (.I0(n2461), .I1(n911), .O(\u_VsyHsyGenerator/pCnt_valueNext[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3807.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3808 (.I0(n2461), .I1(n909), .O(\u_VsyHsyGenerator/pCnt_valueNext[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3808.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3809 (.I0(n2461), .I1(n907), .O(\u_VsyHsyGenerator/pCnt_valueNext[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3809.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3810 (.I0(n2461), .I1(n905), .O(\u_VsyHsyGenerator/pCnt_valueNext[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3810.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3811 (.I0(n2461), .I1(n903), .O(\u_VsyHsyGenerator/pCnt_valueNext[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3811.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3812 (.I0(n2461), .I1(n901), .O(\u_VsyHsyGenerator/pCnt_valueNext[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3812.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3813 (.I0(n2461), .I1(n900), .O(\u_VsyHsyGenerator/pCnt_valueNext[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3813.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3814 (.I0(n1429), .I1(n2496), .I2(n898), .O(\u_VsyHsyGenerator/frameCnt_valueNext[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__3814.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__3815 (.I0(n1429), .I1(n2496), .I2(n896), .O(\u_VsyHsyGenerator/frameCnt_valueNext[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__3815.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__3816 (.I0(n1429), .I1(n2496), .I2(n894), .O(\u_VsyHsyGenerator/frameCnt_valueNext[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__3816.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__3817 (.I0(n1429), .I1(n2496), .I2(n892), .O(\u_VsyHsyGenerator/frameCnt_valueNext[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__3817.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__3818 (.I0(n1429), .I1(n2496), .I2(n890), .O(\u_VsyHsyGenerator/frameCnt_valueNext[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__3818.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__3819 (.I0(n1429), .I1(n2496), .I2(n888), .O(\u_VsyHsyGenerator/frameCnt_valueNext[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__3819.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__3820 (.I0(n1429), .I1(n2496), .I2(n869), .O(\u_VsyHsyGenerator/frameCnt_valueNext[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__3820.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__3821 (.I0(n1429), .I1(n2496), .I2(n766), .O(\u_VsyHsyGenerator/frameCnt_valueNext[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__3821.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__3822 (.I0(n1429), .I1(n2496), .I2(n728), .O(\u_VsyHsyGenerator/frameCnt_valueNext[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__3822.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__3823 (.I0(n1429), .I1(\u_VsyHsyGenerator/vsynDl[0] ), 
            .I2(n2456), .O(\u_VsyHsyGenerator/n681 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hefef */ ;
    defparam LUT__3823.LUTMASK = 16'hefef;
    EFX_LUT4 LUT__3824 (.I0(\u_VsyHsyGenerator/n519 ), .I1(\u_VsyHsyGenerator/hsynDl[0] ), 
            .O(\u_VsyHsyGenerator/n416 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3824.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3825 (.I0(\u_VsyHsyGenerator/n519 ), .I1(\u_VsyHsyGenerator/hsynDl[1] ), 
            .O(\u_VsyHsyGenerator/n415 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3825.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3826 (.I0(\u_VsyHsyGenerator/n519 ), .I1(\u_VsyHsyGenerator/hsynDl[2] ), 
            .O(\u_VsyHsyGenerator/n414 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3826.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3827 (.I0(n1429), .I1(n948), .O(\u_VsyHsyGenerator/hsynCnt_valueNext[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3827.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3828 (.I0(n1429), .I1(n946), .O(\u_VsyHsyGenerator/hsynCnt_valueNext[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3828.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3829 (.I0(n1429), .I1(n930), .O(\u_VsyHsyGenerator/hsynCnt_valueNext[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3829.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3830 (.I0(n1429), .I1(n928), .O(\u_VsyHsyGenerator/hsynCnt_valueNext[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3830.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3831 (.I0(n1429), .I1(n926), .O(\u_VsyHsyGenerator/hsynCnt_valueNext[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3831.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3832 (.I0(n1429), .I1(n924), .O(\u_VsyHsyGenerator/hsynCnt_valueNext[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3832.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3833 (.I0(n1429), .I1(n922), .O(\u_VsyHsyGenerator/hsynCnt_valueNext[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3833.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3834 (.I0(n1429), .I1(n920), .O(\u_VsyHsyGenerator/hsynCnt_valueNext[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3834.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3835 (.I0(n1429), .I1(n919), .O(\u_VsyHsyGenerator/hsynCnt_valueNext[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3835.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3836 (.I0(\u_axi4_ctrl/wframe_index[1] ), .I1(\u_axi4_ctrl/wframe_index[0] ), 
            .O(\u_axi4_ctrl/n323 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3836.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3837 (.I0(\u_axi4_ctrl/wframe_vsync_dly[2] ), .I1(\u_axi4_ctrl/wframe_vsync_dly[3] ), 
            .O(\u_axi4_ctrl/equal_37/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3837.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3838 (.I0(\u_lcd_driver/vcnt[0] ), .I1(\u_lcd_driver/vcnt[1] ), 
            .I2(\u_lcd_driver/vcnt[2] ), .I3(\u_lcd_driver/vcnt[3] ), .O(n2497)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0007 */ ;
    defparam LUT__3838.LUTMASK = 16'h0007;
    EFX_LUT4 LUT__3839 (.I0(\u_lcd_driver/vcnt[4] ), .I1(n2497), .I2(n2441), 
            .O(n2498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3839.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3840 (.I0(\u_lcd_driver/vcnt[5] ), .I1(n2438), .I2(n2498), 
            .O(\u_lcd_driver/n108 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3840.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3841 (.I0(\u_axi4_ctrl/wfifo_cnt[4] ), .I1(\u_axi4_ctrl/wfifo_cnt[3] ), 
            .I2(\u_axi4_ctrl/wfifo_cnt[2] ), .I3(\u_axi4_ctrl/wfifo_cnt[1] ), 
            .O(n2499)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3841.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3842 (.I0(\u_axi4_ctrl/wfifo_cnt[0] ), .I1(n2499), .O(\u_axi4_ctrl/equal_28/n9 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3842.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3843 (.I0(\u_axi4_ctrl/equal_28/n9 ), .I1(n516), .O(\u_axi4_ctrl/n96 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3843.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3844 (.I0(\u_axi4_ctrl/wframe_vsync_dly[3] ), .I1(\u_axi4_ctrl/wframe_vsync_dly[2] ), 
            .I2(\Axi0ResetReg[2] ), .O(\u_axi4_ctrl/n1476 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__3844.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__3845 (.I0(\u_axi4_ctrl/wframe_index[1] ), .I1(\u_axi4_ctrl/wframe_index[0] ), 
            .O(\u_axi4_ctrl/n324 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3845.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3846 (.I0(\u_VsyHsyGenerator/pCnt_value[4] ), .I1(\u_VsyHsyGenerator/pCnt_value[7] ), 
            .I2(\u_VsyHsyGenerator/pCnt_value[9] ), .I3(\u_VsyHsyGenerator/pCnt_value[8] ), 
            .O(n2500)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe7f */ ;
    defparam LUT__3846.LUTMASK = 16'hfe7f;
    EFX_LUT4 LUT__3847 (.I0(\u_VsyHsyGenerator/pCnt_value[9] ), .I1(\u_VsyHsyGenerator/pCnt_value[7] ), 
            .I2(\u_VsyHsyGenerator/pCnt_value[8] ), .I3(\u_VsyHsyGenerator/pCnt_value[4] ), 
            .O(n2501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__3847.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__3848 (.I0(n2501), .I1(n2500), .I2(\u_VsyHsyGenerator/pCnt_value[3] ), 
            .I3(\u_VsyHsyGenerator/pCnt_value[6] ), .O(n2502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf5cf */ ;
    defparam LUT__3848.LUTMASK = 16'hf5cf;
    EFX_LUT4 LUT__3849 (.I0(n2502), .I1(n2480), .I2(\u_VsyHsyGenerator/pCnt_value[5] ), 
            .O(n2503)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3849.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3850 (.I0(n2487), .I1(n2503), .I2(n2481), .I3(n2477), 
            .O(\XYCrop_frame_Gray[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__3850.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__3851 (.I0(\u_axi4_ctrl/wframe_index[0] ), .I1(\u_axi4_ctrl/wframe_index[1] ), 
            .O(\u_axi4_ctrl/n343 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3851.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3852 (.I0(\u_axi4_ctrl/rframe_vsync_dly[2] ), .I1(\u_axi4_ctrl/rframe_vsync_dly[3] ), 
            .O(\u_axi4_ctrl/equal_46/n3 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3852.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3853 (.I0(n2430), .I1(\u_axi4_ctrl/n370 ), .O(n2504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3853.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3854 (.I0(DdrCtrl_BVALID_0), .I1(\u_axi4_ctrl/state[0] ), 
            .I2(\u_axi4_ctrl/state[1] ), .O(n2505)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__3854.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__3855 (.I0(n2504), .I1(n2433), .I2(\u_axi4_ctrl/n1531 ), 
            .I3(n2505), .O(n2506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f00 */ ;
    defparam LUT__3855.LUTMASK = 16'h7f00;
    EFX_LUT4 LUT__3856 (.I0(n257), .I1(n259), .O(n2507)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3856.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3857 (.I0(n261), .I1(n263), .I2(n265), .I3(n761), 
            .O(n2508)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3857.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3858 (.I0(n2508), .I1(n2507), .I2(n255), .I3(n254), 
            .O(n2509)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h008f */ ;
    defparam LUT__3858.LUTMASK = 16'h008f;
    EFX_LUT4 LUT__3859 (.I0(\u_axi4_ctrl/state[0] ), .I1(\u_axi4_ctrl/state[1] ), 
            .I2(\u_axi4_ctrl/state[2] ), .O(n2510)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__3859.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__3860 (.I0(n298), .I1(n300), .I2(n297), .I3(n2510), 
            .O(\u_axi4_ctrl/n412 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfe00 */ ;
    defparam LUT__3860.LUTMASK = 16'hfe00;
    EFX_LUT4 LUT__3861 (.I0(DdrCtrl_AREADY_0), .I1(\u_axi4_ctrl/state[0] ), 
            .I2(\u_axi4_ctrl/state[1] ), .O(n2511)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__3861.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__3862 (.I0(\u_axi4_ctrl/n412 ), .I1(n2509), .I2(n2511), 
            .O(n2512)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hd0d0 */ ;
    defparam LUT__3862.LUTMASK = 16'hd0d0;
    EFX_LUT4 LUT__3863 (.I0(\u_axi4_ctrl/rdata_cnt_dly[6] ), .I1(\u_axi4_ctrl/rdata_cnt_dly[7] ), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[8] ), .O(n2513)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0101 */ ;
    defparam LUT__3863.LUTMASK = 16'h0101;
    EFX_LUT4 LUT__3864 (.I0(\u_axi4_ctrl/rdata_cnt_dly[1] ), .I1(\u_axi4_ctrl/rdata_cnt_dly[0] ), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[2] ), .I3(\u_axi4_ctrl/rdata_cnt_dly[3] ), 
            .O(n2514)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3864.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3865 (.I0(\u_axi4_ctrl/rdata_cnt_dly[4] ), .I1(\u_axi4_ctrl/rdata_cnt_dly[5] ), 
            .O(n2515)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3865.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3866 (.I0(\u_axi4_ctrl/state[1] ), .I1(\u_axi4_ctrl/state[0] ), 
            .I2(DdrCtrl_RVALID_0), .I3(\u_axi4_ctrl/state[2] ), .O(\u_axi4_ctrl/n386 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__3866.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__3867 (.I0(n2513), .I1(n2514), .I2(n2515), .I3(\u_axi4_ctrl/n386 ), 
            .O(\u_axi4_ctrl/n388 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3867.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3868 (.I0(DdrCtrl_AREADY_0), .I1(\u_axi4_ctrl/state[0] ), 
            .I2(\u_axi4_ctrl/n388 ), .I3(n2435), .O(n2516)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e00 */ ;
    defparam LUT__3868.LUTMASK = 16'h0e00;
    EFX_LUT4 LUT__3869 (.I0(n2512), .I1(\u_axi4_ctrl/state[2] ), .I2(n2506), 
            .I3(n2516), .O(\u_axi4_ctrl/n396 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hff01 */ ;
    defparam LUT__3869.LUTMASK = 16'hff01;
    EFX_LUT4 LUT__3870 (.I0(n2509), .I1(n2510), .O(n2517)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3870.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3871 (.I0(n2517), .I1(\Axi0ResetReg[2] ), .O(\u_axi4_ctrl/n1483 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3871.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3872 (.I0(n2474), .I1(n2476), .I2(\u_VsyHsyGenerator/hsynCnt_value[9] ), 
            .O(n2518)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3e3e */ ;
    defparam LUT__3872.LUTMASK = 16'h3e3e;
    EFX_LUT4 LUT__3873 (.I0(\u_VsyHsyGenerator/pCnt_value[3] ), .I1(\u_VsyHsyGenerator/pCnt_value[4] ), 
            .I2(n2462), .I3(n2457), .O(n2519)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__3873.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__3874 (.I0(n2482), .I1(n2519), .I2(n2486), .O(n2520)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3874.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3875 (.I0(n2503), .I1(n2518), .I2(n2484), .I3(n2520), 
            .O(\XYCrop_frame_Gray[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hfeff */ ;
    defparam LUT__3875.LUTMASK = 16'hfeff;
    EFX_LUT4 LUT__3876 (.I0(n2518), .I1(n2520), .O(\XYCrop_frame_Gray[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3876.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3877 (.I0(\u_axi4_ctrl/equal_28/n9 ), .I1(n723), .O(\u_axi4_ctrl/n92 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3877.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3878 (.I0(\u_axi4_ctrl/equal_28/n9 ), .I1(n724), .O(\u_axi4_ctrl/n93 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3878.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3879 (.I0(\u_axi4_ctrl/rdata_cnt_dly[1] ), .I1(\u_axi4_ctrl/rdata_cnt_dly[0] ), 
            .O(\u_axi4_ctrl/n1551 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3879.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3880 (.I0(\u_axi4_ctrl/equal_28/n9 ), .I1(n726), .O(\u_axi4_ctrl/n94 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3880.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3881 (.I0(\u_axi4_ctrl/equal_28/n9 ), .I1(n399), .O(\u_axi4_ctrl/n95 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3881.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3882 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[3] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] ), .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[7] ), 
            .O(n2521)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3882.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3883 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[5] ), 
            .I2(n2521), .O(n2522)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__3883.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__3884 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[0] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] ), .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] ), 
            .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[4] ), 
            .O(n2523)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3884.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3885 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[2] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[11] ), 
            .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[8] ), 
            .O(n2524)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3885.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3886 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[1] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] ), .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.waddr_cntr_sync_g2b_r[6] ), 
            .O(n2525)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3886.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3887 (.I0(n2522), .I1(n2523), .I2(n2524), .I3(n2525), 
            .O(n2526)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3887.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3888 (.I0(lvds_tx2_DATA[0]), .I1(\u_axi4_ctrl/rfifo_empty ), 
            .I2(n2526), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/rd_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0e0e */ ;
    defparam LUT__3888.LUTMASK = 16'h0e0e;
    EFX_LUT4 LUT__3889 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[3] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] ), .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[8] ), 
            .O(n2527)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3889.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3890 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[4] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] ), .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[9] ), 
            .O(n2528)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3890.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3891 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[5] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
            .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[11] ), 
            .O(n2529)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0990 */ ;
    defparam LUT__3891.LUTMASK = 16'h0990;
    EFX_LUT4 LUT__3892 (.I0(n2527), .I1(n2528), .I2(n2529), .O(n2530)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3892.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3893 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[6] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] ), .I3(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[10] ), 
            .O(n2531)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9009 */ ;
    defparam LUT__3893.LUTMASK = 16'h9009;
    EFX_LUT4 LUT__3894 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.genblk1.raddr_cntr_sync_g2b_r[7] ), 
            .I2(n2531), .O(n2532)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9090 */ ;
    defparam LUT__3894.LUTMASK = 16'h9090;
    EFX_LUT4 LUT__3895 (.I0(n2532), .I1(n2530), .I2(\u_axi4_ctrl/rfifo_wenb ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/wr_en_int )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7070 */ ;
    defparam LUT__3895.LUTMASK = 16'h7070;
    EFX_LUT4 LUT__3896 (.I0(n2472), .I1(\u_axi4_ctrl/wfifo_empty ), .I2(\u_axi4_ctrl/n370 ), 
            .O(ceg_net12)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__3896.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__3897 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] ), 
            .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__3897.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__3898 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] ), 
            .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] ), 
            .I3(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6996 */ ;
    defparam LUT__3898.LUTMASK = 16'h6996;
    EFX_LUT4 LUT__3899 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[2] ), 
            .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__3899.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__3900 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[0] ), 
            .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__3900.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__3901 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/raddr[0] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[0] ), 
            .I2(\u_axi4_ctrl/wfifo_empty ), .O(n1776)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3901.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3902 (.I0(n1574), .I1(n1776), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3902.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3905 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[2] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[1] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3905.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3906 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3906.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3907 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3907.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3908 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3908.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3909 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3909.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3910 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[10] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11] ), 
            .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__3910.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__3911 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[10] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] ), 
            .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] ), 
            .I3(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6996 */ ;
    defparam LUT__3911.LUTMASK = 16'h6996;
    EFX_LUT4 LUT__3912 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] ), 
            .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__3912.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__3913 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3] ), 
            .I2(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__3913.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__3914 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3914.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3915 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3915.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3916 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[10] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[9] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3916.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3917 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[9] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3917.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3918 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[11] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[12] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3918.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3919 (.I0(n1571), .I1(n1574), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3919.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3920 (.I0(n1568), .I1(n1571), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3920.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3921 (.I0(n1565), .I1(n1568), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3921.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3922 (.I0(n1562), .I1(n1565), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3922.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3923 (.I0(n1559), .I1(n1562), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3923.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3924 (.I0(n1556), .I1(n1559), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3924.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3925 (.I0(n1553), .I1(n1556), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3925.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3926 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[9] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] ), 
            .I2(\u_axi4_ctrl/wfifo_empty ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3926.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3927 (.I0(n1553), .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_w[9] ), 
            .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__3927.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__3928 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[3] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3928.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3929 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[4] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3929.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3930 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[5] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3930.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3931 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[6] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3931.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3932 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[7] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3932.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3933 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[8] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3933.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3934 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[9] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3934.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3935 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[10] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3935.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3936 (.I0(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[12] ), 
            .I1(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/waddr[11] ), .O(\u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3936.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3937 (.I0(n2526), .I1(\u_axi4_ctrl/rfifo_empty ), .I2(lvds_tx2_DATA[0]), 
            .O(ceg_net19)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0b0b */ ;
    defparam LUT__3937.LUTMASK = 16'h0b0b;
    EFX_LUT4 LUT__3938 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__3938.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__3939 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[4] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__3939.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__3940 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[2] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__3940.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__3941 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[0] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__3941.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__3942 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[0] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3942.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3945 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[9] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__3945.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__3946 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[9] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[7] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__3946.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__3947 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[5] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__3947.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__3948 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[3] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9696 */ ;
    defparam LUT__3948.LUTMASK = 16'h9696;
    EFX_LUT4 LUT__3949 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[5] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[4] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3949.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3950 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[7] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[6] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3950.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3951 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[9] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[8] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3951.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3952 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[10] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry_sync[11] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_sync_g2b[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3952.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3953 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[2] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[1] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3953.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3954 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[4] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[3] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3954.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3955 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[5] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3955.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3956 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[7] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry_sync[8] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_sync_g2b[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3956.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3957 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[3] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] ), 
            .O(n2533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__3957.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__3958 (.I0(n2533), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[3] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] ), .I3(\u_axi4_ctrl/rfifo_empty ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3c55 */ ;
    defparam LUT__3958.LUTMASK = 16'h3c55;
    EFX_LUT4 LUT__3959 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[4] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] ), 
            .O(n2534)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__3959.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__3960 (.I0(n2534), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[4] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] ), .I3(\u_axi4_ctrl/rfifo_empty ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3c55 */ ;
    defparam LUT__3960.LUTMASK = 16'h3c55;
    EFX_LUT4 LUT__3961 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[5] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] ), 
            .O(n2535)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__3961.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__3962 (.I0(n2535), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[5] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] ), .I3(\u_axi4_ctrl/rfifo_empty ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3c55 */ ;
    defparam LUT__3962.LUTMASK = 16'h3c55;
    EFX_LUT4 LUT__3963 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] ), 
            .O(n2536)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__3963.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__3964 (.I0(n2536), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[6] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] ), .I3(\u_axi4_ctrl/rfifo_empty ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3c55 */ ;
    defparam LUT__3964.LUTMASK = 16'h3c55;
    EFX_LUT4 LUT__3965 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[7] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] ), 
            .O(n2537)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__3965.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__3966 (.I0(n2537), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[7] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] ), .I3(\u_axi4_ctrl/rfifo_empty ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3c55 */ ;
    defparam LUT__3966.LUTMASK = 16'h3c55;
    EFX_LUT4 LUT__3967 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[8] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] ), 
            .O(n2538)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__3967.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__3968 (.I0(n2538), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[8] ), 
            .I2(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] ), .I3(\u_axi4_ctrl/rfifo_empty ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3c55 */ ;
    defparam LUT__3968.LUTMASK = 16'h3c55;
    EFX_LUT4 LUT__3969 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[10] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[10] ), 
            .I2(\u_axi4_ctrl/rfifo_empty ), .O(n2539)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3969.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3970 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/raddr[9] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[9] ), 
            .I2(\u_axi4_ctrl/rfifo_empty ), .I3(n2539), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hac53 */ ;
    defparam LUT__3970.LUTMASK = 16'hac53;
    EFX_LUT4 LUT__3971 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr[11] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/raddr_cntr_r[11] ), 
            .I2(\u_axi4_ctrl/rfifo_empty ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3971.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3972 (.I0(n2539), .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[11] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.raddr_cntr_gry[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__3972.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__3973 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[1] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3973.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3974 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[2] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3974.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3975 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[3] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3975.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3976 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[4] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3976.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3977 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[5] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3977.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3978 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[6] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] ), .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3978.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3979 (.I0(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/waddr[7] ), 
            .I1(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/waddr_cntr[8] ), 
            .O(\u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/genblk7.waddr_cntr_gry[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3979.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3980 (.I0(\u_axi4_ctrl/wframe_index[1] ), .I1(\u_axi4_ctrl/wframe_index[0] ), 
            .O(\u_axi4_ctrl/n342 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h9999 */ ;
    defparam LUT__3980.LUTMASK = 16'h9999;
    EFX_LUT4 LUT__3981 (.I0(\u_axi4_ctrl/state[2] ), .I1(\u_axi4_ctrl/state[0] ), 
            .O(n2540)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3981.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3982 (.I0(DdrCtrl_AREADY_0), .I1(DdrCtrl_BVALID_0), .I2(n2540), 
            .I3(\u_axi4_ctrl/state[1] ), .O(\u_axi4_ctrl/n1616 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3fa0 */ ;
    defparam LUT__3982.LUTMASK = 16'h3fa0;
    EFX_LUT4 LUT__3983 (.I0(\u_axi4_ctrl/state[2] ), .I1(\Axi0ResetReg[2] ), 
            .O(\u_axi4_ctrl/n1623 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3983.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3984 (.I0(\u_axi4_ctrl/n388 ), .I1(n2435), .I2(n2517), 
            .O(\u_axi4_ctrl/n394 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf4f4 */ ;
    defparam LUT__3984.LUTMASK = 16'hf4f4;
    EFX_LUT4 LUT__3985 (.I0(DdrCtrl_BREADY_0), .I1(DdrCtrl_BVALID_0), .O(\u_axi4_ctrl/n376 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3985.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3986 (.I0(\u_axi4_ctrl/rframe_vsync_dly[3] ), .I1(\u_axi4_ctrl/rframe_vsync_dly[2] ), 
            .I2(\Axi0ResetReg[2] ), .O(\u_axi4_ctrl/n1485 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4f4f */ ;
    defparam LUT__3986.LUTMASK = 16'h4f4f;
    EFX_LUT4 LUT__3987 (.I0(\u_axi4_ctrl/araddr[10] ), .I1(\u_axi4_ctrl/awaddr[10] ), 
            .I2(n2517), .O(\u_axi4_ctrl/n704 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3987.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3988 (.I0(n2517), .I1(\u_axi4_ctrl/n412 ), .I2(\Axi0ResetReg[2] ), 
            .O(ceg_net124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1010 */ ;
    defparam LUT__3988.LUTMASK = 16'h1010;
    EFX_LUT4 LUT__3989 (.I0(\u_axi4_ctrl/araddr[11] ), .I1(\u_axi4_ctrl/awaddr[11] ), 
            .I2(n2517), .O(\u_axi4_ctrl/n703 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3989.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3990 (.I0(\u_axi4_ctrl/araddr[12] ), .I1(\u_axi4_ctrl/awaddr[12] ), 
            .I2(n2517), .O(\u_axi4_ctrl/n702 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3990.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3991 (.I0(\u_axi4_ctrl/araddr[13] ), .I1(\u_axi4_ctrl/awaddr[13] ), 
            .I2(n2517), .O(\u_axi4_ctrl/n701 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3991.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3992 (.I0(\u_axi4_ctrl/araddr[14] ), .I1(\u_axi4_ctrl/awaddr[14] ), 
            .I2(n2517), .O(\u_axi4_ctrl/n700 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3992.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3993 (.I0(\u_axi4_ctrl/araddr[15] ), .I1(\u_axi4_ctrl/awaddr[15] ), 
            .I2(n2517), .O(\u_axi4_ctrl/n699 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3993.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3994 (.I0(\u_axi4_ctrl/araddr[16] ), .I1(\u_axi4_ctrl/awaddr[16] ), 
            .I2(n2517), .O(\u_axi4_ctrl/n698 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3994.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3995 (.I0(\u_axi4_ctrl/araddr[17] ), .I1(\u_axi4_ctrl/awaddr[17] ), 
            .I2(n2517), .O(\u_axi4_ctrl/n697 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3995.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3996 (.I0(\u_axi4_ctrl/araddr[18] ), .I1(\u_axi4_ctrl/awaddr[18] ), 
            .I2(n2517), .O(\u_axi4_ctrl/n696 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3996.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3997 (.I0(\u_axi4_ctrl/araddr[19] ), .I1(\u_axi4_ctrl/awaddr[19] ), 
            .I2(n2517), .O(\u_axi4_ctrl/n695 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3997.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3998 (.I0(\u_axi4_ctrl/araddr[20] ), .I1(\u_axi4_ctrl/awaddr[20] ), 
            .I2(n2517), .O(\u_axi4_ctrl/n694 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3998.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3999 (.I0(\u_axi4_ctrl/araddr[21] ), .I1(\u_axi4_ctrl/awaddr[21] ), 
            .I2(n2517), .O(\u_axi4_ctrl/n693 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3999.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4000 (.I0(\u_axi4_ctrl/araddr[22] ), .I1(\u_axi4_ctrl/awaddr[22] ), 
            .I2(n2517), .O(\u_axi4_ctrl/n692 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4000.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4001 (.I0(\u_axi4_ctrl/araddr[23] ), .I1(\u_axi4_ctrl/awaddr[23] ), 
            .I2(n2517), .O(\u_axi4_ctrl/n691 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4001.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4002 (.I0(\u_axi4_ctrl/rframe_index[0] ), .I1(\u_axi4_ctrl/wframe_index[0] ), 
            .I2(n2517), .O(\u_axi4_ctrl/n690 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4002.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4003 (.I0(\u_axi4_ctrl/rframe_index[1] ), .I1(\u_axi4_ctrl/wframe_index[1] ), 
            .I2(n2517), .O(\u_axi4_ctrl/n689 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__4003.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__4004 (.I0(\u_axi4_ctrl/wdata_cnt_dly[0] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[1] ), 
            .O(\u_axi4_ctrl/n1506 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__4004.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__4005 (.I0(\u_axi4_ctrl/wdata_cnt_dly[0] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[1] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[2] ), .O(\u_axi4_ctrl/n1511 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__4005.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__4006 (.I0(\u_axi4_ctrl/wdata_cnt_dly[0] ), .I1(\u_axi4_ctrl/wdata_cnt_dly[1] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[2] ), .I3(\u_axi4_ctrl/wdata_cnt_dly[3] ), 
            .O(\u_axi4_ctrl/n1516 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__4006.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__4007 (.I0(n2430), .I1(\u_axi4_ctrl/wdata_cnt_dly[4] ), 
            .O(\u_axi4_ctrl/n1521 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__4007.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__4008 (.I0(n2430), .I1(\u_axi4_ctrl/wdata_cnt_dly[4] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[5] ), .O(\u_axi4_ctrl/n1526 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__4008.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__4009 (.I0(n2430), .I1(n2434), .I2(\u_axi4_ctrl/wdata_cnt_dly[6] ), 
            .O(n2541)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__4009.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__4010 (.I0(n2541), .I1(\u_axi4_ctrl/wdata_cnt_dly[7] ), 
            .O(\u_axi4_ctrl/n1536 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__4010.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__4011 (.I0(n2541), .I1(\u_axi4_ctrl/wdata_cnt_dly[7] ), 
            .I2(\u_axi4_ctrl/wdata_cnt_dly[8] ), .O(\u_axi4_ctrl/n1541 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__4011.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__4012 (.I0(\u_axi4_ctrl/rdata_cnt_dly[1] ), .I1(\u_axi4_ctrl/rdata_cnt_dly[0] ), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[2] ), .O(\u_axi4_ctrl/n1556 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__4012.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__4013 (.I0(\u_axi4_ctrl/rdata_cnt_dly[1] ), .I1(\u_axi4_ctrl/rdata_cnt_dly[0] ), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[2] ), .I3(\u_axi4_ctrl/rdata_cnt_dly[3] ), 
            .O(\u_axi4_ctrl/n1561 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__4013.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__4014 (.I0(n2514), .I1(\u_axi4_ctrl/rdata_cnt_dly[4] ), 
            .O(\u_axi4_ctrl/n1566 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__4014.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__4015 (.I0(n2514), .I1(\u_axi4_ctrl/rdata_cnt_dly[4] ), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[5] ), .O(\u_axi4_ctrl/n1571 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__4015.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__4016 (.I0(n2514), .I1(n2515), .O(n2542)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4016.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4017 (.I0(n2542), .I1(\u_axi4_ctrl/rdata_cnt_dly[6] ), 
            .O(\u_axi4_ctrl/n1576 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__4017.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__4018 (.I0(n2542), .I1(\u_axi4_ctrl/rdata_cnt_dly[6] ), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[7] ), .O(\u_axi4_ctrl/n1581 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__4018.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__4019 (.I0(n2542), .I1(\u_axi4_ctrl/rdata_cnt_dly[6] ), 
            .I2(\u_axi4_ctrl/rdata_cnt_dly[7] ), .I3(\u_axi4_ctrl/rdata_cnt_dly[8] ), 
            .O(\u_axi4_ctrl/n1586 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__4019.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__4020 (.I0(\u_lcd_driver/vcnt[3] ), .I1(\u_lcd_driver/vcnt[4] ), 
            .I2(\u_lcd_driver/vcnt[5] ), .I3(\u_lcd_driver/vcnt[6] ), .O(n2543)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__4020.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__4021 (.I0(\u_lcd_driver/vcnt[2] ), .I1(\u_lcd_driver/vcnt[1] ), 
            .I2(n2543), .I3(n2440), .O(n2544)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__4021.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__4022 (.I0(n2544), .I1(\u_lcd_driver/vcnt[9] ), .I2(n2441), 
            .O(n2545)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hb0b0 */ ;
    defparam LUT__4022.LUTMASK = 16'hb0b0;
    EFX_LUT4 LUT__4023 (.I0(\u_lcd_driver/vcnt[0] ), .I1(n2545), .O(\u_lcd_driver/n81 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__4023.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__4024 (.I0(\u_lcd_driver/hcnt[0] ), .I1(\u_lcd_driver/hcnt[1] ), 
            .O(n2546)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4024.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4025 (.I0(\u_lcd_driver/hcnt[2] ), .I1(\u_lcd_driver/hcnt[3] ), 
            .I2(\u_lcd_driver/hcnt[4] ), .I3(\u_lcd_driver/hcnt[5] ), .O(n2547)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__4025.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__4026 (.I0(\u_lcd_driver/hcnt[6] ), .I1(\u_lcd_driver/hcnt[7] ), 
            .O(n2548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__4026.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__4027 (.I0(\u_lcd_driver/hcnt[9] ), .I1(\u_lcd_driver/hcnt[11] ), 
            .I2(\u_lcd_driver/hcnt[10] ), .I3(\u_lcd_driver/hcnt[8] ), .O(n2549)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__4027.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__4028 (.I0(n2546), .I1(n2547), .I2(n2548), .I3(n2549), 
            .O(\u_lcd_driver/equal_15/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__4028.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__4029 (.I0(n2546), .I1(n2547), .I2(n2548), .I3(\u_lcd_driver/hcnt[8] ), 
            .O(n2550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8f00 */ ;
    defparam LUT__4029.LUTMASK = 16'h8f00;
    EFX_LUT4 LUT__4030 (.I0(n2550), .I1(\u_lcd_driver/hcnt[9] ), .I2(\u_lcd_driver/hcnt[10] ), 
            .I3(\u_lcd_driver/hcnt[11] ), .O(n2551)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__4030.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__4031 (.I0(\u_lcd_driver/hcnt[0] ), .I1(n2551), .O(\u_lcd_driver/n34 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__4031.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__4032 (.I0(n2545), .I1(n1137), .O(\u_lcd_driver/n80 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4032.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4033 (.I0(n2545), .I1(n233), .O(\u_lcd_driver/n79 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4033.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4034 (.I0(n2545), .I1(n231), .O(\u_lcd_driver/n78 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4034.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4035 (.I0(n2545), .I1(n229), .O(\u_lcd_driver/n77 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4035.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4036 (.I0(n2545), .I1(n227), .O(\u_lcd_driver/n76 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4036.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4037 (.I0(n2545), .I1(n225), .O(\u_lcd_driver/n75 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4037.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4038 (.I0(n2545), .I1(n223), .O(\u_lcd_driver/n74 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4038.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4039 (.I0(n2545), .I1(n221), .O(\u_lcd_driver/n73 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4039.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4040 (.I0(n2545), .I1(n219), .O(\u_lcd_driver/n72 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4040.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4041 (.I0(n2545), .I1(n217), .O(\u_lcd_driver/n71 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4041.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4042 (.I0(n2545), .I1(n216), .O(\u_lcd_driver/n70 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4042.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4043 (.I0(n2551), .I1(n776), .O(\u_lcd_driver/n33 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4043.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4044 (.I0(n2551), .I1(n252), .O(\u_lcd_driver/n32 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4044.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4045 (.I0(n2551), .I1(n250), .O(\u_lcd_driver/n31 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4045.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4046 (.I0(n2551), .I1(n248), .O(\u_lcd_driver/n30 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4046.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4047 (.I0(n2551), .I1(n246), .O(\u_lcd_driver/n29 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4047.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4048 (.I0(n2551), .I1(n244), .O(\u_lcd_driver/n28 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4048.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4049 (.I0(n2551), .I1(n242), .O(\u_lcd_driver/n27 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4049.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4050 (.I0(n2551), .I1(n240), .O(\u_lcd_driver/n26 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4050.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4051 (.I0(n2551), .I1(n238), .O(\u_lcd_driver/n25 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4051.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4052 (.I0(n2551), .I1(n236), .O(\u_lcd_driver/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4052.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4053 (.I0(n2551), .I1(n235), .O(\u_lcd_driver/n23 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__4053.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__4122 (.I0(\U0_DDR_Reset/u_ddr_reset_sequencer/rstn_dly[1] ), 
            .O(DdrCtrl_CFG_SEQ_RST)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5555, EFX_ATTRIBUTE_INSTANCE__IS_LUT_SOP_INF_INV=TRUE */ ;
    defparam LUT__4122.LUTMASK = 16'h5555;
    EFX_LUT4 LUT__3685 (.I0(\u_axi4_ctrl/state[1] ), .I1(\u_axi4_ctrl/state[0] ), 
            .I2(\u_axi4_ctrl/state[2] ), .O(DdrCtrl_AVALID_0)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__3685.LUTMASK = 16'h1414;
    EFX_GBUFCE CLKBUF__2 (.CE(1'b1), .I(tx_slowclk), .O(\tx_slowclk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__2.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__1 (.CE(1'b1), .I(clk_12M_i), .O(\clk_12M_i~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__1.CE_POLARITY = 1'b1;
    EFX_GBUFCE CLKBUF__0 (.CE(1'b1), .I(Axi_Clk), .O(\Axi_Clk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__0.CE_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i1  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n2556)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/R0_FIFO\R0_FIFO.v(1256)
    defparam \AUX_ADD_CI__u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_axi4_ctrl/u_R0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_41/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i1  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n2555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1263)
    defparam \AUX_ADD_CI__u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_40/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i4  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n2554)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/W0_FIFO\W0_FIFO.v(1261)
    defparam \AUX_ADD_CI__u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_axi4_ctrl/u_W0_FIFO/u_efx_fifo_top/xefx_fifo_ctl/sub_37/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__u_axi4_ctrl/sub_21/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n2553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:\LearningMaterials\FPGA_Competition\VF-T35F324_Board_HDK_Info_V1.51\06_FPGA_Examples_Image\02_AR0135_DVP_DDR3_LVDS_1024600\Source\axi4_ctrl.v(90)
    defparam \AUX_ADD_CI__u_axi4_ctrl/sub_21/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__u_axi4_ctrl/sub_21/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1  (.I0(1'b1), 
            .I1(1'b1), .CI(1'b0), .CO(n2552)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // D:/LearningMaterials/FPGA_Competition/VF-T35F324_Board_HDK_Info_V1.51/06_FPGA_Examples_Image/02_AR0135_DVP_DDR3_LVDS_1024600/Efinity\ip/etx_ddr3_reset_controller\etx_ddr3_reset_controller.v(166)
    defparam \AUX_ADD_CI__U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__U0_DDR_Reset/u_ddr_reset_sequencer/sub_13/add_2/i1 .I1_POLARITY = 1'b1;
    
endmodule

//
// Verific Verilog Description of module EFX_LUT4_e55454b3_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_e55454b3_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_e55454b3_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_e55454b3_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_e55454b3_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_e55454b3_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_e55454b3_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_e55454b3_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_e55454b3_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_e55454b3_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_e55454b3_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_e55454b3_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_e55454b3_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_e55454b3_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_e55454b3_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_e55454b3_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_e55454b3_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_e55454b3_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__1_8_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__1_8_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__1_8_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__1_8_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__1_8_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__1_8_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__1_8_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__1_8_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__1_8_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__1_8_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__1_8_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__1_8_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__1_8_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__16_2_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__1_8_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__1_8_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__16_2_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__1_8_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__16_2_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__16_2_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__16_2_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__16_2_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__16_2_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_e55454b3__16_2_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_e55454b3_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_GBUFCE_e55454b3_0
// module not written out since it is a black box. 
//

