// Generator : SpinalHDL v1.9.3    git head : 029104c77a54c53f1edda327a3bea333f7d65fd9
// Component : VsyHsyGenerator
// Git hash  : 9db8a52bfc668fe3a2234c919a6525e06b49c734

`timescale 1ns/1ps

module VsyHsyGenerator (
  output reg          io_de,
  output     [15:0]   io_color,
  input               io_nextFrame,
  output     [13:0]   ram_addr,
  input      [15:0]   ram_color,
  output     [4:0]    ram_en,
  input               clk,
  input               reset
);

  wire       [15:0]   picture_color_rgb;
  wire       [13:0]   picture_ram_addr;
  wire       [4:0]    picture_ram_en;
  wire       [9:0]    _zz_hCnt_valueNext;
  wire       [0:0]    _zz_hCnt_valueNext_1;
  wire       [9:0]    _zz_pCnt_valueNext;
  wire       [0:0]    _zz_pCnt_valueNext_1;
  reg                 hCnt_willIncrement;
  reg                 hCnt_willClear;
  reg        [9:0]    hCnt_valueNext;
  reg        [9:0]    hCnt_value;
  wire                hCnt_willOverflowIfInc;
  wire                hCnt_willOverflow;
  reg                 pCnt_willIncrement;
  reg                 pCnt_willClear;
  reg        [9:0]    pCnt_valueNext;
  reg        [9:0]    pCnt_value;
  wire                pCnt_willOverflowIfInc;
  wire                pCnt_willOverflow;
  reg                 frameInterval;
  wire                when_MyTopLevel_l25;

  assign _zz_hCnt_valueNext_1 = hCnt_willIncrement;
  assign _zz_hCnt_valueNext = {9'd0, _zz_hCnt_valueNext_1};
  assign _zz_pCnt_valueNext_1 = pCnt_willIncrement;
  assign _zz_pCnt_valueNext = {9'd0, _zz_pCnt_valueNext_1};
  PictureGenerator picture (
    .coordinate_x (pCnt_value[9:0]        ), //i
    .coordinate_y (hCnt_value[9:0]        ), //i
    .color_rgb    (picture_color_rgb[15:0]), //o
    .ram_color    (ram_color[15:0]        ), //i
    .ram_addr     (picture_ram_addr[13:0] ), //o
    .ram_en       (picture_ram_en[4:0]    ), //o
    .clk          (clk                    ), //i
    .reset        (reset                  )  //i
  );
  always @(*) begin
    hCnt_willIncrement = 1'b0;
    if(pCnt_willOverflow) begin
      hCnt_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    hCnt_willClear = 1'b0;
    if(hCnt_willOverflow) begin
      hCnt_willClear = 1'b1;
    end
  end

  assign hCnt_willOverflowIfInc = (hCnt_value == 10'h258);
  assign hCnt_willOverflow = (hCnt_willOverflowIfInc && hCnt_willIncrement);
  always @(*) begin
    if(hCnt_willOverflow) begin
      hCnt_valueNext = 10'h000;
    end else begin
      hCnt_valueNext = (hCnt_value + _zz_hCnt_valueNext);
    end
    if(hCnt_willClear) begin
      hCnt_valueNext = 10'h000;
    end
  end

  always @(*) begin
    pCnt_willIncrement = 1'b0;
    if(when_MyTopLevel_l25) begin
      pCnt_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    pCnt_willClear = 1'b0;
    if(pCnt_willOverflow) begin
      pCnt_willClear = 1'b1;
    end
  end

  assign pCnt_willOverflowIfInc = (pCnt_value == 10'h3ff);
  assign pCnt_willOverflow = (pCnt_willOverflowIfInc && pCnt_willIncrement);
  always @(*) begin
    pCnt_valueNext = (pCnt_value + _zz_pCnt_valueNext);
    if(pCnt_willClear) begin
      pCnt_valueNext = 10'h000;
    end
  end

  always @(*) begin
    io_de = 1'b0;
    if(when_MyTopLevel_l25) begin
      io_de = 1'b1;
    end
  end

  assign when_MyTopLevel_l25 = (! frameInterval);
  assign io_color = picture_color_rgb;
  assign ram_en = picture_ram_en;
  assign ram_addr = picture_ram_addr;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      hCnt_value <= 10'h000;
      pCnt_value <= 10'h000;
      frameInterval <= 1'b1;
    end else begin
      hCnt_value <= hCnt_valueNext;
      pCnt_value <= pCnt_valueNext;
      if(hCnt_willOverflow) begin
        frameInterval <= 1'b1;
      end
      if(frameInterval) begin
        if(io_nextFrame) begin
          frameInterval <= 1'b0;
        end
      end
    end
  end


endmodule

module PictureGenerator (
  input      [9:0]    coordinate_x,
  input      [9:0]    coordinate_y,
  output reg [15:0]   color_rgb,
  input      [15:0]   ram_color,
  output     [13:0]   ram_addr,
  output reg [4:0]    ram_en,
  input               clk,
  input               reset
);

  reg        [9:0]    rAddr_ram_x;
  reg        [9:0]    rAddr_ram_y;
  wire       [4:0]    rAddr_ram_en;
  wire       [13:0]   rAddr_ram_addr;
  wire       [9:0]    _zz_currXDiv;
  wire       [9:0]    _zz_currYDiv;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_1;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_1_1;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_1_2;
  reg        [7:0]    _zz__zz_when_PictureGenerator_l138;
  wire       [6:0]    _zz__zz_when_PictureGenerator_l138_2;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_3;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_4;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_5;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_6;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_7;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_8;
  wire       [11:0]   _zz_when_PictureGenerator_l78_5;
  wire       [11:0]   _zz_when_PictureGenerator_l78_6;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_1_3;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_1_4;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_1_5;
  reg        [7:0]    _zz__zz_when_PictureGenerator_l138_9;
  wire       [6:0]    _zz__zz_when_PictureGenerator_l138_10;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_11;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_12;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_13;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_14;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_15;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_16;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_17;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_1_6;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_1_7;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_1_8;
  reg        [7:0]    _zz__zz_when_PictureGenerator_l138_18;
  wire       [6:0]    _zz__zz_when_PictureGenerator_l138_19;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_20;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_21;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_22;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_23;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_24;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_25;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_26;
  wire       [11:0]   _zz_when_PictureGenerator_l81;
  wire       [11:0]   _zz_when_PictureGenerator_l81_1;
  wire       [11:0]   _zz_when_PictureGenerator_l87_5;
  wire       [11:0]   _zz_when_PictureGenerator_l87_6;
  wire       [11:0]   _zz_when_PictureGenerator_l87_7;
  wire       [11:0]   _zz_when_PictureGenerator_l87_8;
  wire       [11:0]   _zz_when_PictureGenerator_l87_9;
  wire       [11:0]   _zz_when_PictureGenerator_l87_10;
  wire       [2:0]    _zz_when_PictureGenerator_l138_10;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_3_1;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_3_2;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_3_3;
  reg        [7:0]    _zz__zz_when_PictureGenerator_l138_2_1;
  wire       [6:0]    _zz__zz_when_PictureGenerator_l138_2_2;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_2_3;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_2_4;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_2_5;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_2_6;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_2_7;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_2_8;
  wire       [11:0]   _zz_when_PictureGenerator_l78_1_1;
  wire       [11:0]   _zz_when_PictureGenerator_l78_1_2;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_3_4;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_3_5;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_3_6;
  reg        [7:0]    _zz__zz_when_PictureGenerator_l138_2_9;
  wire       [6:0]    _zz__zz_when_PictureGenerator_l138_2_10;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_2_11;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_2_12;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_2_13;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_2_14;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_2_15;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_2_16;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_2_17;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_3_7;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_3_8;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_3_9;
  reg        [7:0]    _zz__zz_when_PictureGenerator_l138_2_18;
  wire       [6:0]    _zz__zz_when_PictureGenerator_l138_2_19;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_2_20;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_2_21;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_2_22;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_2_23;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_2_24;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_2_25;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_2_26;
  wire       [11:0]   _zz_when_PictureGenerator_l81_1_1;
  wire       [11:0]   _zz_when_PictureGenerator_l81_1_2;
  wire       [11:0]   _zz_when_PictureGenerator_l87_1_1;
  wire       [11:0]   _zz_when_PictureGenerator_l87_1_2;
  wire       [11:0]   _zz_when_PictureGenerator_l87_1_3;
  wire       [11:0]   _zz_when_PictureGenerator_l87_1_4;
  wire       [11:0]   _zz_when_PictureGenerator_l87_1_5;
  wire       [11:0]   _zz_when_PictureGenerator_l87_1_6;
  wire       [2:0]    _zz_when_PictureGenerator_l138_1_1;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_5_1;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_5_2;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_5_3;
  reg        [7:0]    _zz__zz_when_PictureGenerator_l138_4_1;
  wire       [6:0]    _zz__zz_when_PictureGenerator_l138_4_2;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_4_3;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_4_4;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_4_5;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_4_6;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_4_7;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_4_8;
  wire       [11:0]   _zz_when_PictureGenerator_l78_2_1;
  wire       [11:0]   _zz_when_PictureGenerator_l78_2_2;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_5_4;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_5_5;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_5_6;
  reg        [7:0]    _zz__zz_when_PictureGenerator_l138_4_9;
  wire       [6:0]    _zz__zz_when_PictureGenerator_l138_4_10;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_4_11;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_4_12;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_4_13;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_4_14;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_4_15;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_4_16;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_4_17;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_5_7;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_5_8;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_5_9;
  reg        [7:0]    _zz__zz_when_PictureGenerator_l138_4_18;
  wire       [6:0]    _zz__zz_when_PictureGenerator_l138_4_19;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_4_20;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_4_21;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_4_22;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_4_23;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_4_24;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_4_25;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_4_26;
  wire       [11:0]   _zz_when_PictureGenerator_l81_2;
  wire       [11:0]   _zz_when_PictureGenerator_l81_2_1;
  wire       [11:0]   _zz_when_PictureGenerator_l87_2_1;
  wire       [11:0]   _zz_when_PictureGenerator_l87_2_2;
  wire       [11:0]   _zz_when_PictureGenerator_l87_2_3;
  wire       [11:0]   _zz_when_PictureGenerator_l87_2_4;
  wire       [11:0]   _zz_when_PictureGenerator_l87_2_5;
  wire       [11:0]   _zz_when_PictureGenerator_l87_2_6;
  wire       [2:0]    _zz_when_PictureGenerator_l138_2_1;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_7_1;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_7_2;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_7_3;
  reg        [7:0]    _zz__zz_when_PictureGenerator_l138_6_1;
  wire       [6:0]    _zz__zz_when_PictureGenerator_l138_6_2;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_6_3;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_6_4;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_6_5;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_6_6;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_6_7;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_6_8;
  wire       [11:0]   _zz_when_PictureGenerator_l78_3_1;
  wire       [11:0]   _zz_when_PictureGenerator_l78_3_2;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_7_4;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_7_5;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_7_6;
  reg        [7:0]    _zz__zz_when_PictureGenerator_l138_6_9;
  wire       [6:0]    _zz__zz_when_PictureGenerator_l138_6_10;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_6_11;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_6_12;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_6_13;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_6_14;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_6_15;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_6_16;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_6_17;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_7_7;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_7_8;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_7_9;
  reg        [7:0]    _zz__zz_when_PictureGenerator_l138_6_18;
  wire       [6:0]    _zz__zz_when_PictureGenerator_l138_6_19;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_6_20;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_6_21;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_6_22;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_6_23;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_6_24;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_6_25;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_6_26;
  wire       [11:0]   _zz_when_PictureGenerator_l81_3;
  wire       [11:0]   _zz_when_PictureGenerator_l81_3_1;
  wire       [11:0]   _zz_when_PictureGenerator_l87_3_1;
  wire       [11:0]   _zz_when_PictureGenerator_l87_3_2;
  wire       [11:0]   _zz_when_PictureGenerator_l87_3_3;
  wire       [11:0]   _zz_when_PictureGenerator_l87_3_4;
  wire       [11:0]   _zz_when_PictureGenerator_l87_3_5;
  wire       [11:0]   _zz_when_PictureGenerator_l87_3_6;
  wire       [2:0]    _zz_when_PictureGenerator_l138_3_1;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_9_1;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_9_2;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_9_3;
  reg        [7:0]    _zz__zz_when_PictureGenerator_l138_8_1;
  wire       [6:0]    _zz__zz_when_PictureGenerator_l138_8_2;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_8_3;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_8_4;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_8_5;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_8_6;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_8_7;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_8_8;
  wire       [11:0]   _zz_when_PictureGenerator_l78_4_1;
  wire       [11:0]   _zz_when_PictureGenerator_l78_4_2;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_9_4;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_9_5;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_9_6;
  reg        [7:0]    _zz__zz_when_PictureGenerator_l138_8_9;
  wire       [6:0]    _zz__zz_when_PictureGenerator_l138_8_10;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_8_11;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_8_12;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_8_13;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_8_14;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_8_15;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_8_16;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_8_17;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_9_7;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_9_8;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_9_9;
  reg        [7:0]    _zz__zz_when_PictureGenerator_l138_8_18;
  wire       [6:0]    _zz__zz_when_PictureGenerator_l138_8_19;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_8_20;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_8_21;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_8_22;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_8_23;
  wire       [11:0]   _zz__zz_when_PictureGenerator_l138_8_24;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_8_25;
  wire       [9:0]    _zz__zz_when_PictureGenerator_l138_8_26;
  wire       [11:0]   _zz_when_PictureGenerator_l81_4;
  wire       [11:0]   _zz_when_PictureGenerator_l81_4_1;
  wire       [11:0]   _zz_when_PictureGenerator_l87_4_1;
  wire       [11:0]   _zz_when_PictureGenerator_l87_4_2;
  wire       [11:0]   _zz_when_PictureGenerator_l87_4_3;
  wire       [11:0]   _zz_when_PictureGenerator_l87_4_4;
  wire       [11:0]   _zz_when_PictureGenerator_l87_4_5;
  wire       [11:0]   _zz_when_PictureGenerator_l87_4_6;
  wire       [2:0]    _zz_when_PictureGenerator_l138_4_1;
  reg        [15:0]   colorInRam;
  wire       [9:0]    currYDiv;
  wire       [9:0]    currXDiv;
  wire       [7:0]    fontVec_0_0;
  wire       [7:0]    fontVec_0_1;
  wire       [7:0]    fontVec_0_2;
  wire       [7:0]    fontVec_0_3;
  wire       [7:0]    fontVec_0_4;
  wire       [7:0]    fontVec_0_5;
  wire       [7:0]    fontVec_0_6;
  wire       [7:0]    fontVec_0_7;
  wire       [7:0]    fontVec_0_8;
  wire       [7:0]    fontVec_0_9;
  wire       [7:0]    fontVec_0_10;
  wire       [7:0]    fontVec_0_11;
  wire       [7:0]    fontVec_0_12;
  wire       [7:0]    fontVec_0_13;
  wire       [7:0]    fontVec_0_14;
  wire       [7:0]    fontVec_0_15;
  wire       [7:0]    fontVec_0_16;
  wire       [7:0]    fontVec_0_17;
  wire       [7:0]    fontVec_0_18;
  wire       [7:0]    fontVec_0_19;
  wire       [7:0]    fontVec_0_20;
  wire       [7:0]    fontVec_0_21;
  wire       [7:0]    fontVec_0_22;
  wire       [7:0]    fontVec_0_23;
  wire       [7:0]    fontVec_0_24;
  wire       [7:0]    fontVec_0_25;
  wire       [7:0]    fontVec_0_26;
  wire       [7:0]    fontVec_0_27;
  wire       [7:0]    fontVec_0_28;
  wire       [7:0]    fontVec_0_29;
  wire       [7:0]    fontVec_0_30;
  wire       [7:0]    fontVec_0_31;
  wire       [7:0]    fontVec_0_32;
  wire       [7:0]    fontVec_0_33;
  wire       [7:0]    fontVec_0_34;
  wire       [7:0]    fontVec_0_35;
  wire       [7:0]    fontVec_0_36;
  wire       [7:0]    fontVec_0_37;
  wire       [7:0]    fontVec_0_38;
  wire       [7:0]    fontVec_0_39;
  wire       [7:0]    fontVec_0_40;
  wire       [7:0]    fontVec_0_41;
  wire       [7:0]    fontVec_0_42;
  wire       [7:0]    fontVec_0_43;
  wire       [7:0]    fontVec_0_44;
  wire       [7:0]    fontVec_0_45;
  wire       [7:0]    fontVec_0_46;
  wire       [7:0]    fontVec_0_47;
  wire       [7:0]    fontVec_0_48;
  wire       [7:0]    fontVec_0_49;
  wire       [7:0]    fontVec_0_50;
  wire       [7:0]    fontVec_0_51;
  wire       [7:0]    fontVec_0_52;
  wire       [7:0]    fontVec_0_53;
  wire       [7:0]    fontVec_0_54;
  wire       [7:0]    fontVec_0_55;
  wire       [7:0]    fontVec_0_56;
  wire       [7:0]    fontVec_0_57;
  wire       [7:0]    fontVec_0_58;
  wire       [7:0]    fontVec_0_59;
  wire       [7:0]    fontVec_0_60;
  wire       [7:0]    fontVec_0_61;
  wire       [7:0]    fontVec_0_62;
  wire       [7:0]    fontVec_0_63;
  wire       [7:0]    fontVec_0_64;
  wire       [7:0]    fontVec_0_65;
  wire       [7:0]    fontVec_0_66;
  wire       [7:0]    fontVec_0_67;
  wire       [7:0]    fontVec_0_68;
  wire       [7:0]    fontVec_0_69;
  wire       [7:0]    fontVec_0_70;
  wire       [7:0]    fontVec_0_71;
  wire       [7:0]    fontVec_1_0;
  wire       [7:0]    fontVec_1_1;
  wire       [7:0]    fontVec_1_2;
  wire       [7:0]    fontVec_1_3;
  wire       [7:0]    fontVec_1_4;
  wire       [7:0]    fontVec_1_5;
  wire       [7:0]    fontVec_1_6;
  wire       [7:0]    fontVec_1_7;
  wire       [7:0]    fontVec_1_8;
  wire       [7:0]    fontVec_1_9;
  wire       [7:0]    fontVec_1_10;
  wire       [7:0]    fontVec_1_11;
  wire       [7:0]    fontVec_1_12;
  wire       [7:0]    fontVec_1_13;
  wire       [7:0]    fontVec_1_14;
  wire       [7:0]    fontVec_1_15;
  wire       [7:0]    fontVec_1_16;
  wire       [7:0]    fontVec_1_17;
  wire       [7:0]    fontVec_1_18;
  wire       [7:0]    fontVec_1_19;
  wire       [7:0]    fontVec_1_20;
  wire       [7:0]    fontVec_1_21;
  wire       [7:0]    fontVec_1_22;
  wire       [7:0]    fontVec_1_23;
  wire       [7:0]    fontVec_1_24;
  wire       [7:0]    fontVec_1_25;
  wire       [7:0]    fontVec_1_26;
  wire       [7:0]    fontVec_1_27;
  wire       [7:0]    fontVec_1_28;
  wire       [7:0]    fontVec_1_29;
  wire       [7:0]    fontVec_1_30;
  wire       [7:0]    fontVec_1_31;
  wire       [7:0]    fontVec_1_32;
  wire       [7:0]    fontVec_1_33;
  wire       [7:0]    fontVec_1_34;
  wire       [7:0]    fontVec_1_35;
  wire       [7:0]    fontVec_1_36;
  wire       [7:0]    fontVec_1_37;
  wire       [7:0]    fontVec_1_38;
  wire       [7:0]    fontVec_1_39;
  wire       [7:0]    fontVec_1_40;
  wire       [7:0]    fontVec_1_41;
  wire       [7:0]    fontVec_1_42;
  wire       [7:0]    fontVec_1_43;
  wire       [7:0]    fontVec_1_44;
  wire       [7:0]    fontVec_1_45;
  wire       [7:0]    fontVec_1_46;
  wire       [7:0]    fontVec_1_47;
  wire       [7:0]    fontVec_1_48;
  wire       [7:0]    fontVec_1_49;
  wire       [7:0]    fontVec_1_50;
  wire       [7:0]    fontVec_1_51;
  wire       [7:0]    fontVec_1_52;
  wire       [7:0]    fontVec_1_53;
  wire       [7:0]    fontVec_1_54;
  wire       [7:0]    fontVec_1_55;
  wire       [7:0]    fontVec_1_56;
  wire       [7:0]    fontVec_1_57;
  wire       [7:0]    fontVec_1_58;
  wire       [7:0]    fontVec_1_59;
  wire       [7:0]    fontVec_1_60;
  wire       [7:0]    fontVec_1_61;
  wire       [7:0]    fontVec_1_62;
  wire       [7:0]    fontVec_1_63;
  wire       [7:0]    fontVec_1_64;
  wire       [7:0]    fontVec_1_65;
  wire       [7:0]    fontVec_1_66;
  wire       [7:0]    fontVec_1_67;
  wire       [7:0]    fontVec_1_68;
  wire       [7:0]    fontVec_1_69;
  wire       [7:0]    fontVec_1_70;
  wire       [7:0]    fontVec_1_71;
  wire       [7:0]    fontVec_2_0;
  wire       [7:0]    fontVec_2_1;
  wire       [7:0]    fontVec_2_2;
  wire       [7:0]    fontVec_2_3;
  wire       [7:0]    fontVec_2_4;
  wire       [7:0]    fontVec_2_5;
  wire       [7:0]    fontVec_2_6;
  wire       [7:0]    fontVec_2_7;
  wire       [7:0]    fontVec_2_8;
  wire       [7:0]    fontVec_2_9;
  wire       [7:0]    fontVec_2_10;
  wire       [7:0]    fontVec_2_11;
  wire       [7:0]    fontVec_2_12;
  wire       [7:0]    fontVec_2_13;
  wire       [7:0]    fontVec_2_14;
  wire       [7:0]    fontVec_2_15;
  wire       [7:0]    fontVec_2_16;
  wire       [7:0]    fontVec_2_17;
  wire       [7:0]    fontVec_2_18;
  wire       [7:0]    fontVec_2_19;
  wire       [7:0]    fontVec_2_20;
  wire       [7:0]    fontVec_2_21;
  wire       [7:0]    fontVec_2_22;
  wire       [7:0]    fontVec_2_23;
  wire       [7:0]    fontVec_2_24;
  wire       [7:0]    fontVec_2_25;
  wire       [7:0]    fontVec_2_26;
  wire       [7:0]    fontVec_2_27;
  wire       [7:0]    fontVec_2_28;
  wire       [7:0]    fontVec_2_29;
  wire       [7:0]    fontVec_2_30;
  wire       [7:0]    fontVec_2_31;
  wire       [7:0]    fontVec_2_32;
  wire       [7:0]    fontVec_2_33;
  wire       [7:0]    fontVec_2_34;
  wire       [7:0]    fontVec_2_35;
  wire       [7:0]    fontVec_2_36;
  wire       [7:0]    fontVec_2_37;
  wire       [7:0]    fontVec_2_38;
  wire       [7:0]    fontVec_2_39;
  wire       [7:0]    fontVec_2_40;
  wire       [7:0]    fontVec_2_41;
  wire       [7:0]    fontVec_2_42;
  wire       [7:0]    fontVec_2_43;
  wire       [7:0]    fontVec_2_44;
  wire       [7:0]    fontVec_2_45;
  wire       [7:0]    fontVec_2_46;
  wire       [7:0]    fontVec_2_47;
  wire       [7:0]    fontVec_2_48;
  wire       [7:0]    fontVec_2_49;
  wire       [7:0]    fontVec_2_50;
  wire       [7:0]    fontVec_2_51;
  wire       [7:0]    fontVec_2_52;
  wire       [7:0]    fontVec_2_53;
  wire       [7:0]    fontVec_2_54;
  wire       [7:0]    fontVec_2_55;
  wire       [7:0]    fontVec_2_56;
  wire       [7:0]    fontVec_2_57;
  wire       [7:0]    fontVec_2_58;
  wire       [7:0]    fontVec_2_59;
  wire       [7:0]    fontVec_2_60;
  wire       [7:0]    fontVec_2_61;
  wire       [7:0]    fontVec_2_62;
  wire       [7:0]    fontVec_2_63;
  wire       [7:0]    fontVec_2_64;
  wire       [7:0]    fontVec_2_65;
  wire       [7:0]    fontVec_2_66;
  wire       [7:0]    fontVec_2_67;
  wire       [7:0]    fontVec_2_68;
  wire       [7:0]    fontVec_2_69;
  wire       [7:0]    fontVec_2_70;
  wire       [7:0]    fontVec_2_71;
  wire       [7:0]    fontVec_3_0;
  wire       [7:0]    fontVec_3_1;
  wire       [7:0]    fontVec_3_2;
  wire       [7:0]    fontVec_3_3;
  wire       [7:0]    fontVec_3_4;
  wire       [7:0]    fontVec_3_5;
  wire       [7:0]    fontVec_3_6;
  wire       [7:0]    fontVec_3_7;
  wire       [7:0]    fontVec_3_8;
  wire       [7:0]    fontVec_3_9;
  wire       [7:0]    fontVec_3_10;
  wire       [7:0]    fontVec_3_11;
  wire       [7:0]    fontVec_3_12;
  wire       [7:0]    fontVec_3_13;
  wire       [7:0]    fontVec_3_14;
  wire       [7:0]    fontVec_3_15;
  wire       [7:0]    fontVec_3_16;
  wire       [7:0]    fontVec_3_17;
  wire       [7:0]    fontVec_3_18;
  wire       [7:0]    fontVec_3_19;
  wire       [7:0]    fontVec_3_20;
  wire       [7:0]    fontVec_3_21;
  wire       [7:0]    fontVec_3_22;
  wire       [7:0]    fontVec_3_23;
  wire       [7:0]    fontVec_3_24;
  wire       [7:0]    fontVec_3_25;
  wire       [7:0]    fontVec_3_26;
  wire       [7:0]    fontVec_3_27;
  wire       [7:0]    fontVec_3_28;
  wire       [7:0]    fontVec_3_29;
  wire       [7:0]    fontVec_3_30;
  wire       [7:0]    fontVec_3_31;
  wire       [7:0]    fontVec_3_32;
  wire       [7:0]    fontVec_3_33;
  wire       [7:0]    fontVec_3_34;
  wire       [7:0]    fontVec_3_35;
  wire       [7:0]    fontVec_3_36;
  wire       [7:0]    fontVec_3_37;
  wire       [7:0]    fontVec_3_38;
  wire       [7:0]    fontVec_3_39;
  wire       [7:0]    fontVec_3_40;
  wire       [7:0]    fontVec_3_41;
  wire       [7:0]    fontVec_3_42;
  wire       [7:0]    fontVec_3_43;
  wire       [7:0]    fontVec_3_44;
  wire       [7:0]    fontVec_3_45;
  wire       [7:0]    fontVec_3_46;
  wire       [7:0]    fontVec_3_47;
  wire       [7:0]    fontVec_3_48;
  wire       [7:0]    fontVec_3_49;
  wire       [7:0]    fontVec_3_50;
  wire       [7:0]    fontVec_3_51;
  wire       [7:0]    fontVec_3_52;
  wire       [7:0]    fontVec_3_53;
  wire       [7:0]    fontVec_3_54;
  wire       [7:0]    fontVec_3_55;
  wire       [7:0]    fontVec_3_56;
  wire       [7:0]    fontVec_3_57;
  wire       [7:0]    fontVec_3_58;
  wire       [7:0]    fontVec_3_59;
  wire       [7:0]    fontVec_3_60;
  wire       [7:0]    fontVec_3_61;
  wire       [7:0]    fontVec_3_62;
  wire       [7:0]    fontVec_3_63;
  wire       [7:0]    fontVec_3_64;
  wire       [7:0]    fontVec_3_65;
  wire       [7:0]    fontVec_3_66;
  wire       [7:0]    fontVec_3_67;
  wire       [7:0]    fontVec_3_68;
  wire       [7:0]    fontVec_3_69;
  wire       [7:0]    fontVec_3_70;
  wire       [7:0]    fontVec_3_71;
  wire       [7:0]    fontVec_4_0;
  wire       [7:0]    fontVec_4_1;
  wire       [7:0]    fontVec_4_2;
  wire       [7:0]    fontVec_4_3;
  wire       [7:0]    fontVec_4_4;
  wire       [7:0]    fontVec_4_5;
  wire       [7:0]    fontVec_4_6;
  wire       [7:0]    fontVec_4_7;
  wire       [7:0]    fontVec_4_8;
  wire       [7:0]    fontVec_4_9;
  wire       [7:0]    fontVec_4_10;
  wire       [7:0]    fontVec_4_11;
  wire       [7:0]    fontVec_4_12;
  wire       [7:0]    fontVec_4_13;
  wire       [7:0]    fontVec_4_14;
  wire       [7:0]    fontVec_4_15;
  wire       [7:0]    fontVec_4_16;
  wire       [7:0]    fontVec_4_17;
  wire       [7:0]    fontVec_4_18;
  wire       [7:0]    fontVec_4_19;
  wire       [7:0]    fontVec_4_20;
  wire       [7:0]    fontVec_4_21;
  wire       [7:0]    fontVec_4_22;
  wire       [7:0]    fontVec_4_23;
  wire       [7:0]    fontVec_4_24;
  wire       [7:0]    fontVec_4_25;
  wire       [7:0]    fontVec_4_26;
  wire       [7:0]    fontVec_4_27;
  wire       [7:0]    fontVec_4_28;
  wire       [7:0]    fontVec_4_29;
  wire       [7:0]    fontVec_4_30;
  wire       [7:0]    fontVec_4_31;
  wire       [7:0]    fontVec_4_32;
  wire       [7:0]    fontVec_4_33;
  wire       [7:0]    fontVec_4_34;
  wire       [7:0]    fontVec_4_35;
  wire       [7:0]    fontVec_4_36;
  wire       [7:0]    fontVec_4_37;
  wire       [7:0]    fontVec_4_38;
  wire       [7:0]    fontVec_4_39;
  wire       [7:0]    fontVec_4_40;
  wire       [7:0]    fontVec_4_41;
  wire       [7:0]    fontVec_4_42;
  wire       [7:0]    fontVec_4_43;
  wire       [7:0]    fontVec_4_44;
  wire       [7:0]    fontVec_4_45;
  wire       [7:0]    fontVec_4_46;
  wire       [7:0]    fontVec_4_47;
  wire       [7:0]    fontVec_4_48;
  wire       [7:0]    fontVec_4_49;
  wire       [7:0]    fontVec_4_50;
  wire       [7:0]    fontVec_4_51;
  wire       [7:0]    fontVec_4_52;
  wire       [7:0]    fontVec_4_53;
  wire       [7:0]    fontVec_4_54;
  wire       [7:0]    fontVec_4_55;
  wire       [7:0]    fontVec_4_56;
  wire       [7:0]    fontVec_4_57;
  wire       [7:0]    fontVec_4_58;
  wire       [7:0]    fontVec_4_59;
  wire       [7:0]    fontVec_4_60;
  wire       [7:0]    fontVec_4_61;
  wire       [7:0]    fontVec_4_62;
  wire       [7:0]    fontVec_4_63;
  wire       [7:0]    fontVec_4_64;
  wire       [7:0]    fontVec_4_65;
  wire       [7:0]    fontVec_4_66;
  wire       [7:0]    fontVec_4_67;
  wire       [7:0]    fontVec_4_68;
  wire       [7:0]    fontVec_4_69;
  wire       [7:0]    fontVec_4_70;
  wire       [7:0]    fontVec_4_71;
  wire                when_PictureGenerator_l97;
  wire                when_PictureGenerator_l102;
  wire                when_PictureGenerator_l102_1;
  wire                when_PictureGenerator_l102_2;
  wire                when_PictureGenerator_l102_3;
  wire                when_PictureGenerator_l102_4;
  wire                when_PictureGenerator_l102_5;
  wire                when_PictureGenerator_l102_6;
  wire                when_PictureGenerator_l102_7;
  wire                when_PictureGenerator_l102_8;
  wire                when_PictureGenerator_l102_9;
  wire                when_PictureGenerator_l102_10;
  wire                when_PictureGenerator_l102_11;
  wire                when_PictureGenerator_l102_12;
  wire                when_PictureGenerator_l102_13;
  wire                when_PictureGenerator_l102_14;
  wire                when_PictureGenerator_l102_15;
  wire                when_PictureGenerator_l102_16;
  wire                when_PictureGenerator_l102_17;
  wire                when_PictureGenerator_l102_18;
  wire                when_PictureGenerator_l102_19;
  wire                when_PictureGenerator_l102_20;
  wire                when_PictureGenerator_l102_21;
  wire                when_PictureGenerator_l102_22;
  wire                when_PictureGenerator_l102_23;
  wire                when_PictureGenerator_l102_24;
  wire                when_PictureGenerator_l102_25;
  wire                when_PictureGenerator_l102_26;
  wire                when_PictureGenerator_l102_27;
  wire                when_PictureGenerator_l102_28;
  wire                when_PictureGenerator_l102_29;
  wire                when_PictureGenerator_l102_30;
  wire                when_PictureGenerator_l102_31;
  wire                when_PictureGenerator_l102_32;
  wire                when_PictureGenerator_l102_33;
  wire                when_PictureGenerator_l102_34;
  wire                when_PictureGenerator_l102_35;
  wire                when_PictureGenerator_l102_36;
  wire                when_PictureGenerator_l102_37;
  wire                when_PictureGenerator_l102_38;
  wire                when_PictureGenerator_l102_39;
  wire                when_PictureGenerator_l102_40;
  wire                when_PictureGenerator_l102_41;
  wire                when_PictureGenerator_l102_42;
  wire                when_PictureGenerator_l102_43;
  wire                when_PictureGenerator_l102_44;
  wire                when_PictureGenerator_l102_45;
  wire                when_PictureGenerator_l102_46;
  wire                when_PictureGenerator_l102_47;
  wire                when_PictureGenerator_l102_48;
  wire                when_PictureGenerator_l102_49;
  wire                when_PictureGenerator_l102_50;
  wire                when_PictureGenerator_l102_51;
  wire                when_PictureGenerator_l102_52;
  wire                when_PictureGenerator_l102_53;
  wire                when_PictureGenerator_l102_54;
  wire                when_PictureGenerator_l102_55;
  wire                when_PictureGenerator_l102_56;
  wire                when_PictureGenerator_l102_57;
  wire                when_PictureGenerator_l102_58;
  wire                when_PictureGenerator_l102_59;
  wire                when_PictureGenerator_l102_60;
  wire                when_PictureGenerator_l102_61;
  wire                when_PictureGenerator_l102_62;
  wire                when_PictureGenerator_l102_63;
  wire                when_PictureGenerator_l102_64;
  wire                when_PictureGenerator_l102_65;
  wire                when_PictureGenerator_l102_66;
  wire                when_PictureGenerator_l102_67;
  wire                when_PictureGenerator_l102_68;
  wire                when_PictureGenerator_l102_69;
  wire                when_PictureGenerator_l102_70;
  wire                when_PictureGenerator_l102_71;
  wire                when_PictureGenerator_l102_72;
  wire                when_PictureGenerator_l102_73;
  wire                when_PictureGenerator_l102_74;
  wire                when_PictureGenerator_l102_75;
  wire                when_PictureGenerator_l102_76;
  wire                when_PictureGenerator_l102_77;
  wire                when_PictureGenerator_l102_78;
  wire                when_PictureGenerator_l102_79;
  wire                when_PictureGenerator_l102_80;
  wire                when_PictureGenerator_l102_81;
  wire                when_PictureGenerator_l102_82;
  wire                when_PictureGenerator_l102_83;
  wire                when_PictureGenerator_l102_84;
  wire                when_PictureGenerator_l102_85;
  wire                when_PictureGenerator_l102_86;
  wire                when_PictureGenerator_l102_87;
  wire                when_PictureGenerator_l102_88;
  wire                when_PictureGenerator_l102_89;
  wire                when_PictureGenerator_l102_90;
  wire                when_PictureGenerator_l102_91;
  wire                when_PictureGenerator_l102_92;
  wire                when_PictureGenerator_l102_93;
  wire                when_PictureGenerator_l102_94;
  wire                when_PictureGenerator_l102_95;
  wire                when_PictureGenerator_l102_96;
  wire                when_PictureGenerator_l102_97;
  wire                when_PictureGenerator_l102_98;
  wire                when_PictureGenerator_l102_99;
  wire                when_PictureGenerator_l102_100;
  wire                when_PictureGenerator_l102_101;
  wire                when_PictureGenerator_l102_102;
  wire                when_PictureGenerator_l102_103;
  wire                when_PictureGenerator_l102_104;
  wire                when_PictureGenerator_l102_105;
  wire                when_PictureGenerator_l102_106;
  wire                when_PictureGenerator_l102_107;
  wire                when_PictureGenerator_l102_108;
  wire                when_PictureGenerator_l102_109;
  wire                when_PictureGenerator_l102_110;
  wire                when_PictureGenerator_l102_111;
  wire                when_PictureGenerator_l102_112;
  wire                when_PictureGenerator_l102_113;
  wire                when_PictureGenerator_l102_114;
  wire                when_PictureGenerator_l102_115;
  wire                when_PictureGenerator_l102_116;
  wire                when_PictureGenerator_l102_117;
  wire                when_PictureGenerator_l102_118;
  wire                when_PictureGenerator_l102_119;
  wire                when_PictureGenerator_l102_120;
  wire                when_PictureGenerator_l102_121;
  wire                when_PictureGenerator_l102_122;
  wire                when_PictureGenerator_l102_123;
  wire                when_PictureGenerator_l102_124;
  wire                when_PictureGenerator_l102_125;
  wire                when_PictureGenerator_l102_126;
  wire                when_PictureGenerator_l102_127;
  wire                when_PictureGenerator_l102_128;
  wire                when_PictureGenerator_l102_129;
  wire                when_PictureGenerator_l102_130;
  wire                when_PictureGenerator_l102_131;
  wire                when_PictureGenerator_l102_132;
  wire                when_PictureGenerator_l102_133;
  wire                when_PictureGenerator_l102_134;
  wire                when_PictureGenerator_l102_135;
  wire                when_PictureGenerator_l102_136;
  wire                when_PictureGenerator_l102_137;
  wire                when_PictureGenerator_l102_138;
  wire                when_PictureGenerator_l102_139;
  wire                when_PictureGenerator_l102_140;
  wire                when_PictureGenerator_l102_141;
  wire                when_PictureGenerator_l102_142;
  wire                when_PictureGenerator_l102_143;
  wire                when_PictureGenerator_l102_144;
  wire                when_PictureGenerator_l102_145;
  wire                when_PictureGenerator_l102_146;
  wire                when_PictureGenerator_l102_147;
  wire                when_PictureGenerator_l102_148;
  wire                when_PictureGenerator_l102_149;
  wire                when_PictureGenerator_l102_150;
  wire                when_PictureGenerator_l102_151;
  wire                when_PictureGenerator_l102_152;
  wire                when_PictureGenerator_l102_153;
  wire                when_PictureGenerator_l102_154;
  wire                when_PictureGenerator_l102_155;
  wire                when_PictureGenerator_l102_156;
  wire                when_PictureGenerator_l102_157;
  wire                when_PictureGenerator_l102_158;
  wire                when_PictureGenerator_l102_159;
  wire                when_PictureGenerator_l102_160;
  wire                when_PictureGenerator_l102_161;
  wire                when_PictureGenerator_l102_162;
  wire                when_PictureGenerator_l102_163;
  wire                when_PictureGenerator_l102_164;
  wire                when_PictureGenerator_l102_165;
  wire                when_PictureGenerator_l102_166;
  wire                when_PictureGenerator_l102_167;
  wire                when_PictureGenerator_l102_168;
  wire                when_PictureGenerator_l102_169;
  wire                when_PictureGenerator_l102_170;
  wire                when_PictureGenerator_l102_171;
  wire                when_PictureGenerator_l102_172;
  wire                when_PictureGenerator_l102_173;
  wire                when_PictureGenerator_l102_174;
  wire                when_PictureGenerator_l102_175;
  wire                when_PictureGenerator_l102_176;
  wire                when_PictureGenerator_l102_177;
  wire                when_PictureGenerator_l102_178;
  wire                when_PictureGenerator_l102_179;
  wire                when_PictureGenerator_l102_180;
  wire                when_PictureGenerator_l102_181;
  wire                when_PictureGenerator_l102_182;
  wire                when_PictureGenerator_l102_183;
  wire                when_PictureGenerator_l102_184;
  wire                when_PictureGenerator_l102_185;
  wire                when_PictureGenerator_l102_186;
  wire                when_PictureGenerator_l102_187;
  wire                when_PictureGenerator_l102_188;
  wire                when_PictureGenerator_l102_189;
  wire                when_PictureGenerator_l102_190;
  wire                when_PictureGenerator_l102_191;
  wire                when_PictureGenerator_l102_192;
  wire                when_PictureGenerator_l102_193;
  wire                when_PictureGenerator_l102_194;
  wire                when_PictureGenerator_l102_195;
  wire                when_PictureGenerator_l102_196;
  wire                when_PictureGenerator_l102_197;
  wire                when_PictureGenerator_l102_198;
  wire                when_PictureGenerator_l102_199;
  wire                when_PictureGenerator_l102_200;
  wire                when_PictureGenerator_l102_201;
  wire                when_PictureGenerator_l102_202;
  wire                when_PictureGenerator_l102_203;
  wire                when_PictureGenerator_l102_204;
  wire                when_PictureGenerator_l102_205;
  wire                when_PictureGenerator_l102_206;
  wire                when_PictureGenerator_l102_207;
  wire                when_PictureGenerator_l102_208;
  wire                when_PictureGenerator_l102_209;
  wire                when_PictureGenerator_l102_210;
  wire                when_PictureGenerator_l102_211;
  wire                when_PictureGenerator_l102_212;
  wire                when_PictureGenerator_l102_213;
  wire                when_PictureGenerator_l102_214;
  wire                when_PictureGenerator_l102_215;
  wire                when_PictureGenerator_l102_216;
  wire                when_PictureGenerator_l102_217;
  wire                when_PictureGenerator_l102_218;
  wire                when_PictureGenerator_l102_219;
  wire                when_PictureGenerator_l102_220;
  wire                when_PictureGenerator_l102_221;
  wire                when_PictureGenerator_l102_222;
  wire                when_PictureGenerator_l102_223;
  wire                when_PictureGenerator_l102_224;
  wire                when_PictureGenerator_l102_225;
  wire                when_PictureGenerator_l102_226;
  wire                when_PictureGenerator_l102_227;
  wire                when_PictureGenerator_l102_228;
  wire                when_PictureGenerator_l102_229;
  wire                when_PictureGenerator_l102_230;
  wire                when_PictureGenerator_l102_231;
  wire                when_PictureGenerator_l102_232;
  wire                when_PictureGenerator_l102_233;
  wire                when_PictureGenerator_l102_234;
  wire                when_PictureGenerator_l102_235;
  wire                when_PictureGenerator_l102_236;
  wire                when_PictureGenerator_l102_237;
  wire                when_PictureGenerator_l102_238;
  wire                when_PictureGenerator_l102_239;
  wire                when_PictureGenerator_l102_240;
  wire                when_PictureGenerator_l102_241;
  wire                when_PictureGenerator_l102_242;
  wire                when_PictureGenerator_l102_243;
  wire                when_PictureGenerator_l102_244;
  wire                when_PictureGenerator_l102_245;
  wire                when_PictureGenerator_l102_246;
  wire                when_PictureGenerator_l102_247;
  wire                when_PictureGenerator_l102_248;
  wire                when_PictureGenerator_l102_249;
  wire                when_PictureGenerator_l102_250;
  wire                when_PictureGenerator_l102_251;
  wire                when_PictureGenerator_l102_252;
  wire                when_PictureGenerator_l102_253;
  wire                when_PictureGenerator_l102_254;
  wire                when_PictureGenerator_l102_255;
  wire                when_PictureGenerator_l102_256;
  wire                when_PictureGenerator_l102_257;
  wire                when_PictureGenerator_l102_258;
  wire                when_PictureGenerator_l102_259;
  wire                when_PictureGenerator_l102_260;
  wire                when_PictureGenerator_l102_261;
  wire                when_PictureGenerator_l102_262;
  wire                when_PictureGenerator_l102_263;
  wire                when_PictureGenerator_l102_264;
  wire                when_PictureGenerator_l102_265;
  wire                when_PictureGenerator_l102_266;
  wire                when_PictureGenerator_l102_267;
  wire                when_PictureGenerator_l102_268;
  wire                when_PictureGenerator_l102_269;
  wire                when_PictureGenerator_l102_270;
  wire                when_PictureGenerator_l102_271;
  wire                when_PictureGenerator_l102_272;
  wire                when_PictureGenerator_l102_273;
  wire                when_PictureGenerator_l102_274;
  wire                when_PictureGenerator_l102_275;
  wire                when_PictureGenerator_l102_276;
  wire                when_PictureGenerator_l102_277;
  wire                when_PictureGenerator_l102_278;
  wire                when_PictureGenerator_l102_279;
  wire                when_PictureGenerator_l102_280;
  wire                when_PictureGenerator_l102_281;
  wire                when_PictureGenerator_l102_282;
  wire                when_PictureGenerator_l102_283;
  wire                when_PictureGenerator_l102_284;
  wire                when_PictureGenerator_l102_285;
  wire                when_PictureGenerator_l102_286;
  wire                when_PictureGenerator_l102_287;
  wire                when_PictureGenerator_l102_288;
  wire                when_PictureGenerator_l102_289;
  wire                when_PictureGenerator_l102_290;
  wire                when_PictureGenerator_l102_291;
  wire                when_PictureGenerator_l102_292;
  wire                when_PictureGenerator_l102_293;
  wire                when_PictureGenerator_l102_294;
  wire                when_PictureGenerator_l102_295;
  wire                when_PictureGenerator_l102_296;
  wire                when_PictureGenerator_l102_297;
  wire                when_PictureGenerator_l102_298;
  wire                when_PictureGenerator_l102_299;
  wire                when_PictureGenerator_l102_300;
  wire                when_PictureGenerator_l102_301;
  wire                when_PictureGenerator_l102_302;
  wire                when_PictureGenerator_l102_303;
  wire                when_PictureGenerator_l102_304;
  wire                when_PictureGenerator_l102_305;
  wire                when_PictureGenerator_l102_306;
  wire                when_PictureGenerator_l102_307;
  wire                when_PictureGenerator_l102_308;
  wire                when_PictureGenerator_l102_309;
  wire                when_PictureGenerator_l102_310;
  wire                when_PictureGenerator_l102_311;
  wire                when_PictureGenerator_l102_312;
  wire                when_PictureGenerator_l102_313;
  wire                when_PictureGenerator_l102_314;
  wire                when_PictureGenerator_l102_315;
  wire                when_PictureGenerator_l102_316;
  wire                when_PictureGenerator_l102_317;
  wire                when_PictureGenerator_l102_318;
  wire                when_PictureGenerator_l102_319;
  wire                when_PictureGenerator_l102_320;
  wire                when_PictureGenerator_l102_321;
  wire                when_PictureGenerator_l102_322;
  wire                when_PictureGenerator_l102_323;
  wire                when_PictureGenerator_l102_324;
  wire                when_PictureGenerator_l102_325;
  wire                when_PictureGenerator_l102_326;
  wire                when_PictureGenerator_l102_327;
  wire                when_PictureGenerator_l102_328;
  wire                when_PictureGenerator_l102_329;
  wire                when_PictureGenerator_l102_330;
  wire                when_PictureGenerator_l102_331;
  wire                when_PictureGenerator_l102_332;
  wire                when_PictureGenerator_l102_333;
  wire                when_PictureGenerator_l102_334;
  wire                when_PictureGenerator_l102_335;
  wire                when_PictureGenerator_l102_336;
  wire                when_PictureGenerator_l102_337;
  wire                when_PictureGenerator_l102_338;
  wire                when_PictureGenerator_l102_339;
  wire                when_PictureGenerator_l102_340;
  wire                when_PictureGenerator_l102_341;
  wire                when_PictureGenerator_l102_342;
  wire                when_PictureGenerator_l102_343;
  wire                when_PictureGenerator_l102_344;
  wire                when_PictureGenerator_l102_345;
  wire                when_PictureGenerator_l102_346;
  wire                when_PictureGenerator_l102_347;
  wire                when_PictureGenerator_l102_348;
  wire                when_PictureGenerator_l102_349;
  wire                when_PictureGenerator_l102_350;
  wire                when_PictureGenerator_l102_351;
  wire                when_PictureGenerator_l102_352;
  wire                when_PictureGenerator_l102_353;
  wire                when_PictureGenerator_l102_354;
  wire                when_PictureGenerator_l102_355;
  wire                when_PictureGenerator_l102_356;
  wire                when_PictureGenerator_l102_357;
  wire                when_PictureGenerator_l102_358;
  wire                when_PictureGenerator_l102_359;
  wire                when_PictureGenerator_l102_360;
  wire                when_PictureGenerator_l102_361;
  wire                when_PictureGenerator_l102_362;
  wire                when_PictureGenerator_l102_363;
  wire                when_PictureGenerator_l102_364;
  wire                when_PictureGenerator_l102_365;
  wire                when_PictureGenerator_l102_366;
  wire                when_PictureGenerator_l102_367;
  wire                when_PictureGenerator_l102_368;
  wire                when_PictureGenerator_l102_369;
  wire                when_PictureGenerator_l102_370;
  wire                when_PictureGenerator_l102_371;
  wire                when_PictureGenerator_l102_372;
  wire                when_PictureGenerator_l102_373;
  wire                when_PictureGenerator_l102_374;
  wire                when_PictureGenerator_l102_375;
  wire                when_PictureGenerator_l102_376;
  wire                when_PictureGenerator_l102_377;
  wire                when_PictureGenerator_l102_378;
  wire                when_PictureGenerator_l102_379;
  wire                when_PictureGenerator_l102_380;
  wire                when_PictureGenerator_l102_381;
  wire                when_PictureGenerator_l102_382;
  wire                when_PictureGenerator_l102_383;
  wire                when_PictureGenerator_l102_384;
  wire                when_PictureGenerator_l102_385;
  wire                when_PictureGenerator_l102_386;
  wire                when_PictureGenerator_l102_387;
  wire                when_PictureGenerator_l102_388;
  wire                when_PictureGenerator_l102_389;
  wire                when_PictureGenerator_l102_390;
  wire                when_PictureGenerator_l102_391;
  wire                when_PictureGenerator_l102_392;
  wire                when_PictureGenerator_l102_393;
  wire                when_PictureGenerator_l102_394;
  wire                when_PictureGenerator_l102_395;
  wire                when_PictureGenerator_l102_396;
  wire                when_PictureGenerator_l102_397;
  wire                when_PictureGenerator_l102_398;
  wire                when_PictureGenerator_l102_399;
  wire                when_PictureGenerator_l102_400;
  wire                when_PictureGenerator_l102_401;
  wire                when_PictureGenerator_l102_402;
  wire                when_PictureGenerator_l102_403;
  wire                when_PictureGenerator_l102_404;
  wire                when_PictureGenerator_l102_405;
  wire                when_PictureGenerator_l102_406;
  wire                when_PictureGenerator_l102_407;
  wire                when_PictureGenerator_l102_408;
  wire                when_PictureGenerator_l102_409;
  wire                when_PictureGenerator_l102_410;
  wire                when_PictureGenerator_l102_411;
  wire                when_PictureGenerator_l102_412;
  wire                when_PictureGenerator_l102_413;
  wire                when_PictureGenerator_l102_414;
  wire                when_PictureGenerator_l102_415;
  wire                when_PictureGenerator_l102_416;
  wire                when_PictureGenerator_l102_417;
  wire                when_PictureGenerator_l102_418;
  wire                when_PictureGenerator_l102_419;
  wire                when_PictureGenerator_l102_420;
  wire                when_PictureGenerator_l102_421;
  wire                when_PictureGenerator_l102_422;
  wire                when_PictureGenerator_l102_423;
  wire                when_PictureGenerator_l102_424;
  wire                when_PictureGenerator_l102_425;
  wire                when_PictureGenerator_l102_426;
  wire                when_PictureGenerator_l102_427;
  wire                when_PictureGenerator_l102_428;
  wire                when_PictureGenerator_l102_429;
  wire                when_PictureGenerator_l102_430;
  wire                when_PictureGenerator_l102_431;
  wire                when_PictureGenerator_l102_432;
  wire                when_PictureGenerator_l102_433;
  wire                when_PictureGenerator_l102_434;
  wire                when_PictureGenerator_l102_435;
  wire                when_PictureGenerator_l102_436;
  wire                when_PictureGenerator_l102_437;
  wire                when_PictureGenerator_l102_438;
  wire                when_PictureGenerator_l102_439;
  wire                when_PictureGenerator_l102_440;
  wire                when_PictureGenerator_l102_441;
  wire                when_PictureGenerator_l102_442;
  wire                when_PictureGenerator_l102_443;
  wire                when_PictureGenerator_l102_444;
  wire                when_PictureGenerator_l102_445;
  wire                when_PictureGenerator_l102_446;
  wire                when_PictureGenerator_l102_447;
  wire                when_PictureGenerator_l102_448;
  wire                when_PictureGenerator_l102_449;
  wire                when_PictureGenerator_l102_450;
  wire                when_PictureGenerator_l102_451;
  wire                when_PictureGenerator_l102_452;
  wire                when_PictureGenerator_l102_453;
  wire                when_PictureGenerator_l102_454;
  wire                when_PictureGenerator_l102_455;
  wire                when_PictureGenerator_l102_456;
  wire                when_PictureGenerator_l102_457;
  wire                when_PictureGenerator_l102_458;
  wire                when_PictureGenerator_l102_459;
  wire                when_PictureGenerator_l102_460;
  wire                when_PictureGenerator_l102_461;
  wire                when_PictureGenerator_l102_462;
  wire                when_PictureGenerator_l102_463;
  wire                when_PictureGenerator_l102_464;
  wire                when_PictureGenerator_l102_465;
  wire                when_PictureGenerator_l102_466;
  wire                when_PictureGenerator_l102_467;
  wire                when_PictureGenerator_l102_468;
  wire                when_PictureGenerator_l102_469;
  wire                when_PictureGenerator_l102_470;
  wire                when_PictureGenerator_l102_471;
  wire                when_PictureGenerator_l102_472;
  wire                when_PictureGenerator_l102_473;
  wire                when_PictureGenerator_l102_474;
  wire                when_PictureGenerator_l102_475;
  wire                when_PictureGenerator_l102_476;
  wire                when_PictureGenerator_l102_477;
  wire                when_PictureGenerator_l102_478;
  wire                when_PictureGenerator_l102_479;
  wire                when_PictureGenerator_l102_480;
  wire                when_PictureGenerator_l102_481;
  wire                when_PictureGenerator_l102_482;
  wire                when_PictureGenerator_l102_483;
  wire                when_PictureGenerator_l102_484;
  wire                when_PictureGenerator_l102_485;
  wire                when_PictureGenerator_l102_486;
  wire                when_PictureGenerator_l102_487;
  wire                when_PictureGenerator_l102_488;
  wire                when_PictureGenerator_l102_489;
  wire                when_PictureGenerator_l102_490;
  wire                when_PictureGenerator_l102_491;
  wire                when_PictureGenerator_l102_492;
  wire                when_PictureGenerator_l102_493;
  wire                when_PictureGenerator_l102_494;
  wire                when_PictureGenerator_l102_495;
  wire                when_PictureGenerator_l102_496;
  wire                when_PictureGenerator_l102_497;
  wire                when_PictureGenerator_l102_498;
  wire                when_PictureGenerator_l102_499;
  wire                when_PictureGenerator_l102_500;
  wire                when_PictureGenerator_l102_501;
  wire                when_PictureGenerator_l102_502;
  wire                when_PictureGenerator_l102_503;
  wire                when_PictureGenerator_l102_504;
  wire                when_PictureGenerator_l102_505;
  wire                when_PictureGenerator_l102_506;
  wire                when_PictureGenerator_l102_507;
  wire                when_PictureGenerator_l102_508;
  wire                when_PictureGenerator_l102_509;
  wire                when_PictureGenerator_l102_510;
  wire                when_PictureGenerator_l102_511;
  wire                when_PictureGenerator_l102_512;
  wire                when_PictureGenerator_l102_513;
  wire                when_PictureGenerator_l102_514;
  wire                when_PictureGenerator_l102_515;
  wire                when_PictureGenerator_l102_516;
  wire                when_PictureGenerator_l102_517;
  wire                when_PictureGenerator_l102_518;
  wire                when_PictureGenerator_l102_519;
  wire                when_PictureGenerator_l102_520;
  wire                when_PictureGenerator_l102_521;
  wire                when_PictureGenerator_l102_522;
  wire                when_PictureGenerator_l102_523;
  wire                when_PictureGenerator_l102_524;
  wire                when_PictureGenerator_l102_525;
  wire                when_PictureGenerator_l102_526;
  wire                when_PictureGenerator_l102_527;
  wire                when_PictureGenerator_l102_528;
  wire                when_PictureGenerator_l102_529;
  wire                when_PictureGenerator_l102_530;
  wire                when_PictureGenerator_l102_531;
  wire                when_PictureGenerator_l102_532;
  wire                when_PictureGenerator_l102_533;
  wire                when_PictureGenerator_l102_534;
  wire                when_PictureGenerator_l102_535;
  wire                when_PictureGenerator_l102_536;
  wire                when_PictureGenerator_l102_537;
  wire                when_PictureGenerator_l102_538;
  wire                when_PictureGenerator_l102_539;
  wire                when_PictureGenerator_l102_540;
  wire                when_PictureGenerator_l102_541;
  wire                when_PictureGenerator_l102_542;
  wire                when_PictureGenerator_l102_543;
  wire                when_PictureGenerator_l102_544;
  wire                when_PictureGenerator_l102_545;
  wire                when_PictureGenerator_l102_546;
  wire                when_PictureGenerator_l102_547;
  wire                when_PictureGenerator_l102_548;
  wire                when_PictureGenerator_l102_549;
  wire                when_PictureGenerator_l102_550;
  wire                when_PictureGenerator_l102_551;
  wire                when_PictureGenerator_l102_552;
  wire                when_PictureGenerator_l102_553;
  wire                when_PictureGenerator_l102_554;
  wire                when_PictureGenerator_l102_555;
  wire                when_PictureGenerator_l102_556;
  wire                when_PictureGenerator_l102_557;
  wire                when_PictureGenerator_l102_558;
  wire                when_PictureGenerator_l102_559;
  wire                when_PictureGenerator_l102_560;
  wire                when_PictureGenerator_l102_561;
  wire                when_PictureGenerator_l102_562;
  wire                when_PictureGenerator_l102_563;
  wire                when_PictureGenerator_l102_564;
  wire                when_PictureGenerator_l102_565;
  wire                when_PictureGenerator_l102_566;
  wire                when_PictureGenerator_l102_567;
  wire                when_PictureGenerator_l102_568;
  wire                when_PictureGenerator_l102_569;
  wire                when_PictureGenerator_l102_570;
  wire                when_PictureGenerator_l102_571;
  wire                when_PictureGenerator_l102_572;
  wire                when_PictureGenerator_l102_573;
  wire                when_PictureGenerator_l102_574;
  wire                when_PictureGenerator_l102_575;
  wire                when_PictureGenerator_l102_576;
  wire                when_PictureGenerator_l102_577;
  wire                when_PictureGenerator_l102_578;
  wire                when_PictureGenerator_l102_579;
  wire                when_PictureGenerator_l102_580;
  wire                when_PictureGenerator_l102_581;
  wire                when_PictureGenerator_l102_582;
  wire                when_PictureGenerator_l102_583;
  wire                when_PictureGenerator_l102_584;
  wire                when_PictureGenerator_l102_585;
  wire                when_PictureGenerator_l102_586;
  wire                when_PictureGenerator_l102_587;
  wire                when_PictureGenerator_l102_588;
  wire                when_PictureGenerator_l102_589;
  wire                when_PictureGenerator_l102_590;
  wire                when_PictureGenerator_l102_591;
  wire                when_PictureGenerator_l102_592;
  wire                when_PictureGenerator_l102_593;
  wire                when_PictureGenerator_l102_594;
  wire                when_PictureGenerator_l102_595;
  wire                when_PictureGenerator_l102_596;
  wire                when_PictureGenerator_l102_597;
  wire                when_PictureGenerator_l102_598;
  wire                when_PictureGenerator_l102_599;
  wire                when_PictureGenerator_l102_600;
  wire                when_PictureGenerator_l102_601;
  wire                when_PictureGenerator_l102_602;
  wire                when_PictureGenerator_l102_603;
  wire                when_PictureGenerator_l102_604;
  wire                when_PictureGenerator_l102_605;
  wire                when_PictureGenerator_l102_606;
  wire                when_PictureGenerator_l102_607;
  wire                when_PictureGenerator_l102_608;
  wire                when_PictureGenerator_l102_609;
  wire                when_PictureGenerator_l102_610;
  wire                when_PictureGenerator_l102_611;
  wire                when_PictureGenerator_l102_612;
  wire                when_PictureGenerator_l102_613;
  wire                when_PictureGenerator_l102_614;
  wire                when_PictureGenerator_l102_615;
  wire                when_PictureGenerator_l102_616;
  wire                when_PictureGenerator_l102_617;
  wire                when_PictureGenerator_l102_618;
  wire                when_PictureGenerator_l102_619;
  wire                when_PictureGenerator_l102_620;
  wire                when_PictureGenerator_l102_621;
  wire                when_PictureGenerator_l102_622;
  wire                when_PictureGenerator_l102_623;
  wire                when_PictureGenerator_l102_624;
  wire                when_PictureGenerator_l102_625;
  wire                when_PictureGenerator_l102_626;
  wire                when_PictureGenerator_l102_627;
  wire                when_PictureGenerator_l102_628;
  wire                when_PictureGenerator_l102_629;
  wire                when_PictureGenerator_l110;
  wire                when_PictureGenerator_l110_1;
  wire                when_PictureGenerator_l110_2;
  wire                when_PictureGenerator_l110_3;
  wire                when_PictureGenerator_l110_4;
  wire                when_PictureGenerator_l110_5;
  wire                when_PictureGenerator_l110_6;
  wire                when_PictureGenerator_l110_7;
  wire                when_PictureGenerator_l110_8;
  wire                when_PictureGenerator_l110_9;
  wire                when_PictureGenerator_l110_10;
  wire                when_PictureGenerator_l110_11;
  wire                when_PictureGenerator_l110_12;
  wire                when_PictureGenerator_l110_13;
  wire                when_PictureGenerator_l110_14;
  wire                when_PictureGenerator_l110_15;
  wire                when_PictureGenerator_l110_16;
  wire                when_PictureGenerator_l110_17;
  wire                when_PictureGenerator_l110_18;
  wire                when_PictureGenerator_l110_19;
  wire                when_PictureGenerator_l110_20;
  wire                when_PictureGenerator_l110_21;
  wire                when_PictureGenerator_l110_22;
  wire                when_PictureGenerator_l110_23;
  wire                when_PictureGenerator_l110_24;
  wire                when_PictureGenerator_l110_25;
  wire                when_PictureGenerator_l110_26;
  wire                when_PictureGenerator_l110_27;
  wire                when_PictureGenerator_l110_28;
  wire                when_PictureGenerator_l110_29;
  wire                when_PictureGenerator_l110_30;
  wire                when_PictureGenerator_l110_31;
  wire                when_PictureGenerator_l110_32;
  wire                when_PictureGenerator_l110_33;
  wire                when_PictureGenerator_l110_34;
  wire                when_PictureGenerator_l110_35;
  wire                when_PictureGenerator_l110_36;
  wire                when_PictureGenerator_l110_37;
  wire                when_PictureGenerator_l110_38;
  wire                when_PictureGenerator_l110_39;
  wire                when_PictureGenerator_l110_40;
  wire                when_PictureGenerator_l110_41;
  wire                when_PictureGenerator_l110_42;
  wire                when_PictureGenerator_l110_43;
  wire                when_PictureGenerator_l110_44;
  wire                when_PictureGenerator_l110_45;
  wire                when_PictureGenerator_l110_46;
  wire                when_PictureGenerator_l110_47;
  wire                when_PictureGenerator_l110_48;
  wire                when_PictureGenerator_l110_49;
  wire                when_PictureGenerator_l110_50;
  wire                when_PictureGenerator_l110_51;
  wire                when_PictureGenerator_l110_52;
  wire                when_PictureGenerator_l110_53;
  wire                when_PictureGenerator_l110_54;
  wire                when_PictureGenerator_l110_55;
  wire                when_PictureGenerator_l110_56;
  wire                when_PictureGenerator_l110_57;
  wire                when_PictureGenerator_l110_58;
  wire                when_PictureGenerator_l110_59;
  wire                when_PictureGenerator_l110_60;
  wire                when_PictureGenerator_l110_61;
  wire                when_PictureGenerator_l110_62;
  wire                when_PictureGenerator_l110_63;
  wire                when_PictureGenerator_l110_64;
  wire                when_PictureGenerator_l110_65;
  wire                when_PictureGenerator_l110_66;
  wire                when_PictureGenerator_l110_67;
  wire                when_PictureGenerator_l110_68;
  wire                when_PictureGenerator_l110_69;
  wire                when_PictureGenerator_l110_70;
  wire                when_PictureGenerator_l110_71;
  wire                when_PictureGenerator_l110_72;
  wire                when_PictureGenerator_l110_73;
  wire                when_PictureGenerator_l110_74;
  wire                when_PictureGenerator_l110_75;
  wire                when_PictureGenerator_l110_76;
  wire                when_PictureGenerator_l110_77;
  wire                when_PictureGenerator_l110_78;
  wire                when_PictureGenerator_l110_79;
  wire                when_PictureGenerator_l110_80;
  wire                when_PictureGenerator_l110_81;
  wire                when_PictureGenerator_l110_82;
  wire                when_PictureGenerator_l110_83;
  wire                when_PictureGenerator_l110_84;
  wire                when_PictureGenerator_l110_85;
  wire                when_PictureGenerator_l110_86;
  wire                when_PictureGenerator_l110_87;
  wire                when_PictureGenerator_l110_88;
  wire                when_PictureGenerator_l110_89;
  wire                when_PictureGenerator_l110_90;
  wire                when_PictureGenerator_l110_91;
  wire                when_PictureGenerator_l110_92;
  wire                when_PictureGenerator_l110_93;
  wire                when_PictureGenerator_l110_94;
  wire                when_PictureGenerator_l110_95;
  wire                when_PictureGenerator_l110_96;
  wire                when_PictureGenerator_l110_97;
  wire                when_PictureGenerator_l110_98;
  wire                when_PictureGenerator_l110_99;
  wire                when_PictureGenerator_l110_100;
  wire                when_PictureGenerator_l110_101;
  wire                when_PictureGenerator_l110_102;
  wire                when_PictureGenerator_l110_103;
  wire                when_PictureGenerator_l110_104;
  wire                when_PictureGenerator_l110_105;
  wire                when_PictureGenerator_l110_106;
  wire                when_PictureGenerator_l110_107;
  wire                when_PictureGenerator_l110_108;
  wire                when_PictureGenerator_l110_109;
  wire                when_PictureGenerator_l110_110;
  wire                when_PictureGenerator_l110_111;
  wire                when_PictureGenerator_l110_112;
  wire                when_PictureGenerator_l110_113;
  wire                when_PictureGenerator_l110_114;
  wire                when_PictureGenerator_l110_115;
  wire                when_PictureGenerator_l110_116;
  wire                when_PictureGenerator_l110_117;
  wire                when_PictureGenerator_l110_118;
  wire                when_PictureGenerator_l110_119;
  wire                when_PictureGenerator_l110_120;
  wire                when_PictureGenerator_l110_121;
  wire                when_PictureGenerator_l110_122;
  wire                when_PictureGenerator_l110_123;
  wire                when_PictureGenerator_l110_124;
  wire                when_PictureGenerator_l110_125;
  wire                when_PictureGenerator_l110_126;
  wire                when_PictureGenerator_l110_127;
  wire                when_PictureGenerator_l110_128;
  wire                when_PictureGenerator_l110_129;
  wire                when_PictureGenerator_l110_130;
  wire                when_PictureGenerator_l110_131;
  wire                when_PictureGenerator_l110_132;
  wire                when_PictureGenerator_l110_133;
  wire                when_PictureGenerator_l110_134;
  wire                when_PictureGenerator_l110_135;
  wire                when_PictureGenerator_l110_136;
  wire                when_PictureGenerator_l110_137;
  wire                when_PictureGenerator_l110_138;
  wire                when_PictureGenerator_l110_139;
  wire                when_PictureGenerator_l110_140;
  wire                when_PictureGenerator_l110_141;
  wire                when_PictureGenerator_l110_142;
  wire                when_PictureGenerator_l110_143;
  wire                when_PictureGenerator_l110_144;
  wire                when_PictureGenerator_l110_145;
  wire                when_PictureGenerator_l110_146;
  wire                when_PictureGenerator_l110_147;
  wire                when_PictureGenerator_l110_148;
  wire                when_PictureGenerator_l110_149;
  wire                when_PictureGenerator_l110_150;
  wire                when_PictureGenerator_l110_151;
  wire                when_PictureGenerator_l110_152;
  wire                when_PictureGenerator_l110_153;
  wire                when_PictureGenerator_l110_154;
  wire                when_PictureGenerator_l110_155;
  wire                when_PictureGenerator_l110_156;
  wire                when_PictureGenerator_l110_157;
  wire                when_PictureGenerator_l110_158;
  wire                when_PictureGenerator_l110_159;
  wire                when_PictureGenerator_l110_160;
  wire                when_PictureGenerator_l110_161;
  wire                when_PictureGenerator_l110_162;
  wire                when_PictureGenerator_l110_163;
  wire                when_PictureGenerator_l110_164;
  wire                when_PictureGenerator_l110_165;
  wire                when_PictureGenerator_l110_166;
  wire                when_PictureGenerator_l110_167;
  wire                when_PictureGenerator_l110_168;
  wire                when_PictureGenerator_l110_169;
  wire                when_PictureGenerator_l110_170;
  wire                when_PictureGenerator_l110_171;
  wire                when_PictureGenerator_l110_172;
  wire                when_PictureGenerator_l110_173;
  wire                when_PictureGenerator_l110_174;
  wire                when_PictureGenerator_l110_175;
  wire                when_PictureGenerator_l110_176;
  wire                when_PictureGenerator_l110_177;
  wire                when_PictureGenerator_l110_178;
  wire                when_PictureGenerator_l110_179;
  wire                when_PictureGenerator_l110_180;
  wire                when_PictureGenerator_l110_181;
  wire                when_PictureGenerator_l110_182;
  wire                when_PictureGenerator_l110_183;
  wire                when_PictureGenerator_l110_184;
  wire                when_PictureGenerator_l110_185;
  wire                when_PictureGenerator_l110_186;
  wire                when_PictureGenerator_l110_187;
  wire                when_PictureGenerator_l110_188;
  wire                when_PictureGenerator_l110_189;
  wire                when_PictureGenerator_l110_190;
  wire                when_PictureGenerator_l110_191;
  wire                when_PictureGenerator_l110_192;
  wire                when_PictureGenerator_l110_193;
  wire                when_PictureGenerator_l110_194;
  wire                when_PictureGenerator_l110_195;
  wire                when_PictureGenerator_l110_196;
  wire                when_PictureGenerator_l110_197;
  wire                when_PictureGenerator_l110_198;
  wire                when_PictureGenerator_l110_199;
  wire                when_PictureGenerator_l110_200;
  wire                when_PictureGenerator_l110_201;
  wire                when_PictureGenerator_l110_202;
  wire                when_PictureGenerator_l110_203;
  wire                when_PictureGenerator_l110_204;
  wire                when_PictureGenerator_l110_205;
  wire                when_PictureGenerator_l110_206;
  wire                when_PictureGenerator_l110_207;
  wire                when_PictureGenerator_l110_208;
  wire                when_PictureGenerator_l110_209;
  wire                when_PictureGenerator_l110_210;
  wire                when_PictureGenerator_l110_211;
  wire                when_PictureGenerator_l110_212;
  wire                when_PictureGenerator_l110_213;
  wire                when_PictureGenerator_l110_214;
  wire                when_PictureGenerator_l110_215;
  wire                when_PictureGenerator_l110_216;
  wire                when_PictureGenerator_l110_217;
  wire                when_PictureGenerator_l110_218;
  wire                when_PictureGenerator_l110_219;
  wire                when_PictureGenerator_l110_220;
  wire                when_PictureGenerator_l110_221;
  wire                when_PictureGenerator_l110_222;
  wire                when_PictureGenerator_l110_223;
  wire                when_PictureGenerator_l110_224;
  wire                when_PictureGenerator_l110_225;
  wire                when_PictureGenerator_l110_226;
  wire                when_PictureGenerator_l110_227;
  wire                when_PictureGenerator_l110_228;
  wire                when_PictureGenerator_l110_229;
  wire                when_PictureGenerator_l110_230;
  wire                when_PictureGenerator_l110_231;
  wire                when_PictureGenerator_l110_232;
  wire                when_PictureGenerator_l110_233;
  wire                when_PictureGenerator_l110_234;
  wire                when_PictureGenerator_l110_235;
  wire                when_PictureGenerator_l110_236;
  wire                when_PictureGenerator_l110_237;
  wire                when_PictureGenerator_l110_238;
  wire                when_PictureGenerator_l110_239;
  wire                when_PictureGenerator_l110_240;
  wire                when_PictureGenerator_l110_241;
  wire                when_PictureGenerator_l110_242;
  wire                when_PictureGenerator_l110_243;
  wire                when_PictureGenerator_l110_244;
  wire                when_PictureGenerator_l110_245;
  wire                when_PictureGenerator_l110_246;
  wire                when_PictureGenerator_l110_247;
  wire                when_PictureGenerator_l110_248;
  wire                when_PictureGenerator_l110_249;
  wire                when_PictureGenerator_l110_250;
  wire                when_PictureGenerator_l110_251;
  wire                when_PictureGenerator_l110_252;
  wire                when_PictureGenerator_l110_253;
  wire                when_PictureGenerator_l110_254;
  wire                when_PictureGenerator_l110_255;
  wire                when_PictureGenerator_l110_256;
  wire                when_PictureGenerator_l110_257;
  wire                when_PictureGenerator_l110_258;
  wire                when_PictureGenerator_l110_259;
  wire                when_PictureGenerator_l110_260;
  wire                when_PictureGenerator_l110_261;
  wire                when_PictureGenerator_l110_262;
  wire                when_PictureGenerator_l110_263;
  wire                when_PictureGenerator_l110_264;
  wire                when_PictureGenerator_l110_265;
  wire                when_PictureGenerator_l110_266;
  wire                when_PictureGenerator_l110_267;
  wire                when_PictureGenerator_l110_268;
  wire                when_PictureGenerator_l110_269;
  wire                when_PictureGenerator_l110_270;
  wire                when_PictureGenerator_l110_271;
  wire                when_PictureGenerator_l110_272;
  wire                when_PictureGenerator_l110_273;
  wire                when_PictureGenerator_l110_274;
  wire                when_PictureGenerator_l110_275;
  wire                when_PictureGenerator_l110_276;
  wire                when_PictureGenerator_l110_277;
  wire                when_PictureGenerator_l110_278;
  wire                when_PictureGenerator_l110_279;
  wire                when_PictureGenerator_l110_280;
  wire                when_PictureGenerator_l110_281;
  wire                when_PictureGenerator_l110_282;
  wire                when_PictureGenerator_l110_283;
  wire                when_PictureGenerator_l110_284;
  wire                when_PictureGenerator_l110_285;
  wire                when_PictureGenerator_l110_286;
  wire                when_PictureGenerator_l110_287;
  wire                when_PictureGenerator_l110_288;
  wire                when_PictureGenerator_l110_289;
  wire                when_PictureGenerator_l110_290;
  wire                when_PictureGenerator_l110_291;
  wire                when_PictureGenerator_l110_292;
  wire                when_PictureGenerator_l110_293;
  wire                when_PictureGenerator_l110_294;
  wire                when_PictureGenerator_l110_295;
  wire                when_PictureGenerator_l110_296;
  wire                when_PictureGenerator_l110_297;
  wire                when_PictureGenerator_l110_298;
  wire                when_PictureGenerator_l110_299;
  wire                when_PictureGenerator_l110_300;
  wire                when_PictureGenerator_l110_301;
  wire                when_PictureGenerator_l110_302;
  wire                when_PictureGenerator_l110_303;
  wire                when_PictureGenerator_l110_304;
  wire                when_PictureGenerator_l110_305;
  wire                when_PictureGenerator_l110_306;
  wire                when_PictureGenerator_l110_307;
  wire                when_PictureGenerator_l110_308;
  wire                when_PictureGenerator_l110_309;
  wire                when_PictureGenerator_l110_310;
  wire                when_PictureGenerator_l110_311;
  wire                when_PictureGenerator_l110_312;
  wire                when_PictureGenerator_l110_313;
  wire                when_PictureGenerator_l110_314;
  wire                when_PictureGenerator_l110_315;
  wire                when_PictureGenerator_l110_316;
  wire                when_PictureGenerator_l110_317;
  wire                when_PictureGenerator_l110_318;
  wire                when_PictureGenerator_l110_319;
  wire                when_PictureGenerator_l110_320;
  wire                when_PictureGenerator_l110_321;
  wire                when_PictureGenerator_l110_322;
  wire                when_PictureGenerator_l110_323;
  wire                when_PictureGenerator_l110_324;
  wire                when_PictureGenerator_l110_325;
  wire                when_PictureGenerator_l110_326;
  wire                when_PictureGenerator_l110_327;
  wire                when_PictureGenerator_l110_328;
  wire                when_PictureGenerator_l110_329;
  wire                when_PictureGenerator_l110_330;
  wire                when_PictureGenerator_l110_331;
  wire                when_PictureGenerator_l110_332;
  wire                when_PictureGenerator_l110_333;
  wire                when_PictureGenerator_l110_334;
  wire                when_PictureGenerator_l110_335;
  wire                when_PictureGenerator_l110_336;
  wire                when_PictureGenerator_l110_337;
  wire                when_PictureGenerator_l110_338;
  wire                when_PictureGenerator_l110_339;
  wire                when_PictureGenerator_l110_340;
  wire                when_PictureGenerator_l110_341;
  wire                when_PictureGenerator_l110_342;
  wire                when_PictureGenerator_l110_343;
  wire                when_PictureGenerator_l110_344;
  wire                when_PictureGenerator_l110_345;
  wire                when_PictureGenerator_l110_346;
  wire                when_PictureGenerator_l110_347;
  wire                when_PictureGenerator_l110_348;
  wire                when_PictureGenerator_l110_349;
  wire                when_PictureGenerator_l110_350;
  wire                when_PictureGenerator_l110_351;
  wire                when_PictureGenerator_l110_352;
  wire                when_PictureGenerator_l110_353;
  wire                when_PictureGenerator_l110_354;
  wire                when_PictureGenerator_l110_355;
  wire                when_PictureGenerator_l110_356;
  wire                when_PictureGenerator_l110_357;
  wire                when_PictureGenerator_l110_358;
  wire                when_PictureGenerator_l110_359;
  wire                when_PictureGenerator_l110_360;
  wire                when_PictureGenerator_l110_361;
  wire                when_PictureGenerator_l110_362;
  wire                when_PictureGenerator_l110_363;
  wire                when_PictureGenerator_l110_364;
  wire                when_PictureGenerator_l110_365;
  wire                when_PictureGenerator_l110_366;
  wire                when_PictureGenerator_l110_367;
  wire                when_PictureGenerator_l110_368;
  wire                when_PictureGenerator_l110_369;
  wire                when_PictureGenerator_l110_370;
  wire                when_PictureGenerator_l110_371;
  wire                when_PictureGenerator_l110_372;
  wire                when_PictureGenerator_l110_373;
  wire                when_PictureGenerator_l110_374;
  wire                when_PictureGenerator_l110_375;
  wire                when_PictureGenerator_l110_376;
  wire                when_PictureGenerator_l110_377;
  wire                when_PictureGenerator_l110_378;
  wire                when_PictureGenerator_l110_379;
  wire                when_PictureGenerator_l110_380;
  wire                when_PictureGenerator_l110_381;
  wire                when_PictureGenerator_l110_382;
  wire                when_PictureGenerator_l110_383;
  wire                when_PictureGenerator_l110_384;
  wire                when_PictureGenerator_l110_385;
  wire                when_PictureGenerator_l110_386;
  wire                when_PictureGenerator_l110_387;
  wire                when_PictureGenerator_l110_388;
  wire                when_PictureGenerator_l110_389;
  wire                when_PictureGenerator_l110_390;
  wire                when_PictureGenerator_l110_391;
  wire                when_PictureGenerator_l110_392;
  wire                when_PictureGenerator_l110_393;
  wire                when_PictureGenerator_l110_394;
  wire                when_PictureGenerator_l110_395;
  wire                when_PictureGenerator_l110_396;
  wire                when_PictureGenerator_l110_397;
  wire                when_PictureGenerator_l110_398;
  wire                when_PictureGenerator_l110_399;
  wire                when_PictureGenerator_l110_400;
  wire                when_PictureGenerator_l110_401;
  wire                when_PictureGenerator_l110_402;
  wire                when_PictureGenerator_l110_403;
  wire                when_PictureGenerator_l110_404;
  wire                when_PictureGenerator_l110_405;
  wire                when_PictureGenerator_l110_406;
  wire                when_PictureGenerator_l110_407;
  wire                when_PictureGenerator_l110_408;
  wire                when_PictureGenerator_l110_409;
  wire                when_PictureGenerator_l110_410;
  wire                when_PictureGenerator_l110_411;
  wire                when_PictureGenerator_l110_412;
  wire                when_PictureGenerator_l110_413;
  wire                when_PictureGenerator_l110_414;
  wire                when_PictureGenerator_l110_415;
  wire                when_PictureGenerator_l110_416;
  wire                when_PictureGenerator_l110_417;
  wire                when_PictureGenerator_l110_418;
  wire                when_PictureGenerator_l110_419;
  wire                when_PictureGenerator_l110_420;
  wire                when_PictureGenerator_l110_421;
  wire                when_PictureGenerator_l110_422;
  wire                when_PictureGenerator_l110_423;
  wire                when_PictureGenerator_l110_424;
  wire                when_PictureGenerator_l110_425;
  wire                when_PictureGenerator_l110_426;
  wire                when_PictureGenerator_l110_427;
  wire                when_PictureGenerator_l110_428;
  wire                when_PictureGenerator_l110_429;
  wire                when_PictureGenerator_l110_430;
  wire                when_PictureGenerator_l110_431;
  wire                when_PictureGenerator_l110_432;
  wire                when_PictureGenerator_l110_433;
  wire                when_PictureGenerator_l110_434;
  wire                when_PictureGenerator_l110_435;
  wire                when_PictureGenerator_l110_436;
  wire                when_PictureGenerator_l110_437;
  wire                when_PictureGenerator_l110_438;
  wire                when_PictureGenerator_l110_439;
  wire                when_PictureGenerator_l110_440;
  wire                when_PictureGenerator_l110_441;
  wire                when_PictureGenerator_l110_442;
  wire                when_PictureGenerator_l110_443;
  wire                when_PictureGenerator_l110_444;
  wire                when_PictureGenerator_l110_445;
  wire                when_PictureGenerator_l110_446;
  wire                when_PictureGenerator_l110_447;
  wire                when_PictureGenerator_l110_448;
  wire                when_PictureGenerator_l110_449;
  wire                when_PictureGenerator_l110_450;
  wire                when_PictureGenerator_l110_451;
  wire                when_PictureGenerator_l110_452;
  wire                when_PictureGenerator_l110_453;
  wire                when_PictureGenerator_l110_454;
  wire                when_PictureGenerator_l110_455;
  wire                when_PictureGenerator_l110_456;
  wire                when_PictureGenerator_l110_457;
  wire                when_PictureGenerator_l110_458;
  wire                when_PictureGenerator_l110_459;
  wire                when_PictureGenerator_l110_460;
  wire                when_PictureGenerator_l110_461;
  wire                when_PictureGenerator_l110_462;
  wire                when_PictureGenerator_l110_463;
  wire                when_PictureGenerator_l110_464;
  wire                when_PictureGenerator_l110_465;
  wire                when_PictureGenerator_l110_466;
  wire                when_PictureGenerator_l110_467;
  wire                when_PictureGenerator_l110_468;
  wire                when_PictureGenerator_l110_469;
  wire                when_PictureGenerator_l110_470;
  wire                when_PictureGenerator_l110_471;
  wire                when_PictureGenerator_l110_472;
  wire                when_PictureGenerator_l110_473;
  wire                when_PictureGenerator_l110_474;
  wire                when_PictureGenerator_l110_475;
  wire                when_PictureGenerator_l110_476;
  wire                when_PictureGenerator_l110_477;
  wire                when_PictureGenerator_l110_478;
  wire                when_PictureGenerator_l110_479;
  wire                when_PictureGenerator_l110_480;
  wire                when_PictureGenerator_l110_481;
  wire                when_PictureGenerator_l110_482;
  wire                when_PictureGenerator_l110_483;
  wire                when_PictureGenerator_l110_484;
  wire                when_PictureGenerator_l110_485;
  wire                when_PictureGenerator_l110_486;
  wire                when_PictureGenerator_l110_487;
  wire                when_PictureGenerator_l110_488;
  wire                when_PictureGenerator_l110_489;
  wire                when_PictureGenerator_l110_490;
  wire                when_PictureGenerator_l110_491;
  wire                when_PictureGenerator_l110_492;
  wire                when_PictureGenerator_l110_493;
  wire                when_PictureGenerator_l110_494;
  wire                when_PictureGenerator_l110_495;
  wire                when_PictureGenerator_l110_496;
  wire                when_PictureGenerator_l110_497;
  wire                when_PictureGenerator_l110_498;
  wire                when_PictureGenerator_l110_499;
  wire                when_PictureGenerator_l110_500;
  wire                when_PictureGenerator_l110_501;
  wire                when_PictureGenerator_l110_502;
  wire                when_PictureGenerator_l110_503;
  wire                when_PictureGenerator_l110_504;
  wire                when_PictureGenerator_l110_505;
  wire                when_PictureGenerator_l110_506;
  wire                when_PictureGenerator_l110_507;
  wire                when_PictureGenerator_l110_508;
  wire                when_PictureGenerator_l110_509;
  wire                when_PictureGenerator_l110_510;
  wire                when_PictureGenerator_l110_511;
  wire                when_PictureGenerator_l110_512;
  wire                when_PictureGenerator_l110_513;
  wire                when_PictureGenerator_l110_514;
  wire                when_PictureGenerator_l110_515;
  wire                when_PictureGenerator_l110_516;
  wire                when_PictureGenerator_l110_517;
  wire                when_PictureGenerator_l115;
  wire                when_PictureGenerator_l117;
  wire                when_PictureGenerator_l119;
  wire                when_PictureGenerator_l121;
  wire                when_PictureGenerator_l130;
  reg        [7:0]    _zz_when_PictureGenerator_l138;
  reg        [7:0]    _zz_when_PictureGenerator_l138_1;
  wire       [11:0]   _zz_when_PictureGenerator_l78;
  wire       [11:0]   _zz_when_PictureGenerator_l87;
  reg                 when_PictureGenerator_l138;
  wire                when_PictureGenerator_l78;
  wire                when_PictureGenerator_l81;
  wire                when_PictureGenerator_l87;
  reg        [7:0]    _zz_when_PictureGenerator_l138_2;
  reg        [7:0]    _zz_when_PictureGenerator_l138_3;
  wire       [11:0]   _zz_when_PictureGenerator_l78_1;
  wire       [11:0]   _zz_when_PictureGenerator_l87_1;
  reg                 when_PictureGenerator_l138_1;
  wire                when_PictureGenerator_l78_1;
  wire                when_PictureGenerator_l81_1;
  wire                when_PictureGenerator_l87_1;
  reg        [7:0]    _zz_when_PictureGenerator_l138_4;
  reg        [7:0]    _zz_when_PictureGenerator_l138_5;
  wire       [11:0]   _zz_when_PictureGenerator_l78_2;
  wire       [11:0]   _zz_when_PictureGenerator_l87_2;
  reg                 when_PictureGenerator_l138_2;
  wire                when_PictureGenerator_l78_2;
  wire                when_PictureGenerator_l81_2;
  wire                when_PictureGenerator_l87_2;
  reg        [7:0]    _zz_when_PictureGenerator_l138_6;
  reg        [7:0]    _zz_when_PictureGenerator_l138_7;
  wire       [11:0]   _zz_when_PictureGenerator_l78_3;
  wire       [11:0]   _zz_when_PictureGenerator_l87_3;
  reg                 when_PictureGenerator_l138_3;
  wire                when_PictureGenerator_l78_3;
  wire                when_PictureGenerator_l81_3;
  wire                when_PictureGenerator_l87_3;
  reg        [7:0]    _zz_when_PictureGenerator_l138_8;
  reg        [7:0]    _zz_when_PictureGenerator_l138_9;
  wire       [11:0]   _zz_when_PictureGenerator_l78_4;
  wire       [11:0]   _zz_when_PictureGenerator_l87_4;
  reg                 when_PictureGenerator_l138_4;
  wire                when_PictureGenerator_l78_4;
  wire                when_PictureGenerator_l81_4;
  wire                when_PictureGenerator_l87_4;

  assign _zz_currXDiv = (coordinate_x >>> 1);
  assign _zz_currYDiv = (coordinate_y >>> 1);
  assign _zz__zz_when_PictureGenerator_l138_1 = (_zz__zz_when_PictureGenerator_l138_1_1 + _zz_when_PictureGenerator_l78);
  assign _zz__zz_when_PictureGenerator_l138_1_2 = (10'h007 - coordinate_x);
  assign _zz__zz_when_PictureGenerator_l138_1_1 = {2'd0, _zz__zz_when_PictureGenerator_l138_1_2};
  assign _zz__zz_when_PictureGenerator_l138_3 = (_zz__zz_when_PictureGenerator_l138_4 - _zz_when_PictureGenerator_l87);
  assign _zz__zz_when_PictureGenerator_l138_2 = _zz__zz_when_PictureGenerator_l138_3[6:0];
  assign _zz__zz_when_PictureGenerator_l138_4 = (_zz__zz_when_PictureGenerator_l138_5 - _zz_when_PictureGenerator_l87);
  assign _zz__zz_when_PictureGenerator_l138_5 = (_zz__zz_when_PictureGenerator_l138_6 - _zz_when_PictureGenerator_l87);
  assign _zz__zz_when_PictureGenerator_l138_7 = (_zz__zz_when_PictureGenerator_l138_8 + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_6 = {2'd0, _zz__zz_when_PictureGenerator_l138_7};
  assign _zz__zz_when_PictureGenerator_l138_8 = (coordinate_y + coordinate_y);
  assign _zz_when_PictureGenerator_l78_5 = (_zz_when_PictureGenerator_l78 + 12'h00f);
  assign _zz_when_PictureGenerator_l78_6 = {2'd0, coordinate_x};
  assign _zz__zz_when_PictureGenerator_l138_1_3 = (_zz__zz_when_PictureGenerator_l138_1_4 + _zz_when_PictureGenerator_l78);
  assign _zz__zz_when_PictureGenerator_l138_1_5 = (10'h017 - coordinate_x);
  assign _zz__zz_when_PictureGenerator_l138_1_4 = {2'd0, _zz__zz_when_PictureGenerator_l138_1_5};
  assign _zz__zz_when_PictureGenerator_l138_11 = (12'h002 + _zz__zz_when_PictureGenerator_l138_12);
  assign _zz__zz_when_PictureGenerator_l138_10 = _zz__zz_when_PictureGenerator_l138_11[6:0];
  assign _zz__zz_when_PictureGenerator_l138_12 = (_zz__zz_when_PictureGenerator_l138_13 - _zz_when_PictureGenerator_l87);
  assign _zz__zz_when_PictureGenerator_l138_13 = (_zz__zz_when_PictureGenerator_l138_14 - _zz_when_PictureGenerator_l87);
  assign _zz__zz_when_PictureGenerator_l138_14 = (_zz__zz_when_PictureGenerator_l138_15 - _zz_when_PictureGenerator_l87);
  assign _zz__zz_when_PictureGenerator_l138_16 = (_zz__zz_when_PictureGenerator_l138_17 + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_15 = {2'd0, _zz__zz_when_PictureGenerator_l138_16};
  assign _zz__zz_when_PictureGenerator_l138_17 = (coordinate_y + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_1_6 = (_zz__zz_when_PictureGenerator_l138_1_7 + _zz_when_PictureGenerator_l78);
  assign _zz__zz_when_PictureGenerator_l138_1_8 = (10'h00f - coordinate_x);
  assign _zz__zz_when_PictureGenerator_l138_1_7 = {2'd0, _zz__zz_when_PictureGenerator_l138_1_8};
  assign _zz__zz_when_PictureGenerator_l138_20 = (12'h001 + _zz__zz_when_PictureGenerator_l138_21);
  assign _zz__zz_when_PictureGenerator_l138_19 = _zz__zz_when_PictureGenerator_l138_20[6:0];
  assign _zz__zz_when_PictureGenerator_l138_21 = (_zz__zz_when_PictureGenerator_l138_22 - _zz_when_PictureGenerator_l87);
  assign _zz__zz_when_PictureGenerator_l138_22 = (_zz__zz_when_PictureGenerator_l138_23 - _zz_when_PictureGenerator_l87);
  assign _zz__zz_when_PictureGenerator_l138_23 = (_zz__zz_when_PictureGenerator_l138_24 - _zz_when_PictureGenerator_l87);
  assign _zz__zz_when_PictureGenerator_l138_25 = (_zz__zz_when_PictureGenerator_l138_26 + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_24 = {2'd0, _zz__zz_when_PictureGenerator_l138_25};
  assign _zz__zz_when_PictureGenerator_l138_26 = (coordinate_y + coordinate_y);
  assign _zz_when_PictureGenerator_l81 = (_zz_when_PictureGenerator_l78 + 12'h007);
  assign _zz_when_PictureGenerator_l81_1 = {2'd0, coordinate_x};
  assign _zz_when_PictureGenerator_l87_5 = {2'd0, coordinate_x};
  assign _zz_when_PictureGenerator_l87_6 = {2'd0, coordinate_y};
  assign _zz_when_PictureGenerator_l87_7 = {2'd0, coordinate_x};
  assign _zz_when_PictureGenerator_l87_8 = (_zz_when_PictureGenerator_l78 + 12'h018);
  assign _zz_when_PictureGenerator_l87_9 = {2'd0, coordinate_y};
  assign _zz_when_PictureGenerator_l87_10 = (_zz_when_PictureGenerator_l87 + 12'h018);
  assign _zz_when_PictureGenerator_l138_10 = _zz_when_PictureGenerator_l138_1[2:0];
  assign _zz__zz_when_PictureGenerator_l138_3_1 = (_zz__zz_when_PictureGenerator_l138_3_2 + _zz_when_PictureGenerator_l78_1);
  assign _zz__zz_when_PictureGenerator_l138_3_3 = (10'h007 - coordinate_x);
  assign _zz__zz_when_PictureGenerator_l138_3_2 = {2'd0, _zz__zz_when_PictureGenerator_l138_3_3};
  assign _zz__zz_when_PictureGenerator_l138_2_3 = (_zz__zz_when_PictureGenerator_l138_2_4 - _zz_when_PictureGenerator_l87_1);
  assign _zz__zz_when_PictureGenerator_l138_2_2 = _zz__zz_when_PictureGenerator_l138_2_3[6:0];
  assign _zz__zz_when_PictureGenerator_l138_2_4 = (_zz__zz_when_PictureGenerator_l138_2_5 - _zz_when_PictureGenerator_l87_1);
  assign _zz__zz_when_PictureGenerator_l138_2_5 = (_zz__zz_when_PictureGenerator_l138_2_6 - _zz_when_PictureGenerator_l87_1);
  assign _zz__zz_when_PictureGenerator_l138_2_7 = (_zz__zz_when_PictureGenerator_l138_2_8 + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_2_6 = {2'd0, _zz__zz_when_PictureGenerator_l138_2_7};
  assign _zz__zz_when_PictureGenerator_l138_2_8 = (coordinate_y + coordinate_y);
  assign _zz_when_PictureGenerator_l78_1_1 = (_zz_when_PictureGenerator_l78_1 + 12'h00f);
  assign _zz_when_PictureGenerator_l78_1_2 = {2'd0, coordinate_x};
  assign _zz__zz_when_PictureGenerator_l138_3_4 = (_zz__zz_when_PictureGenerator_l138_3_5 + _zz_when_PictureGenerator_l78_1);
  assign _zz__zz_when_PictureGenerator_l138_3_6 = (10'h017 - coordinate_x);
  assign _zz__zz_when_PictureGenerator_l138_3_5 = {2'd0, _zz__zz_when_PictureGenerator_l138_3_6};
  assign _zz__zz_when_PictureGenerator_l138_2_11 = (12'h002 + _zz__zz_when_PictureGenerator_l138_2_12);
  assign _zz__zz_when_PictureGenerator_l138_2_10 = _zz__zz_when_PictureGenerator_l138_2_11[6:0];
  assign _zz__zz_when_PictureGenerator_l138_2_12 = (_zz__zz_when_PictureGenerator_l138_2_13 - _zz_when_PictureGenerator_l87_1);
  assign _zz__zz_when_PictureGenerator_l138_2_13 = (_zz__zz_when_PictureGenerator_l138_2_14 - _zz_when_PictureGenerator_l87_1);
  assign _zz__zz_when_PictureGenerator_l138_2_14 = (_zz__zz_when_PictureGenerator_l138_2_15 - _zz_when_PictureGenerator_l87_1);
  assign _zz__zz_when_PictureGenerator_l138_2_16 = (_zz__zz_when_PictureGenerator_l138_2_17 + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_2_15 = {2'd0, _zz__zz_when_PictureGenerator_l138_2_16};
  assign _zz__zz_when_PictureGenerator_l138_2_17 = (coordinate_y + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_3_7 = (_zz__zz_when_PictureGenerator_l138_3_8 + _zz_when_PictureGenerator_l78_1);
  assign _zz__zz_when_PictureGenerator_l138_3_9 = (10'h00f - coordinate_x);
  assign _zz__zz_when_PictureGenerator_l138_3_8 = {2'd0, _zz__zz_when_PictureGenerator_l138_3_9};
  assign _zz__zz_when_PictureGenerator_l138_2_20 = (12'h001 + _zz__zz_when_PictureGenerator_l138_2_21);
  assign _zz__zz_when_PictureGenerator_l138_2_19 = _zz__zz_when_PictureGenerator_l138_2_20[6:0];
  assign _zz__zz_when_PictureGenerator_l138_2_21 = (_zz__zz_when_PictureGenerator_l138_2_22 - _zz_when_PictureGenerator_l87_1);
  assign _zz__zz_when_PictureGenerator_l138_2_22 = (_zz__zz_when_PictureGenerator_l138_2_23 - _zz_when_PictureGenerator_l87_1);
  assign _zz__zz_when_PictureGenerator_l138_2_23 = (_zz__zz_when_PictureGenerator_l138_2_24 - _zz_when_PictureGenerator_l87_1);
  assign _zz__zz_when_PictureGenerator_l138_2_25 = (_zz__zz_when_PictureGenerator_l138_2_26 + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_2_24 = {2'd0, _zz__zz_when_PictureGenerator_l138_2_25};
  assign _zz__zz_when_PictureGenerator_l138_2_26 = (coordinate_y + coordinate_y);
  assign _zz_when_PictureGenerator_l81_1_1 = (_zz_when_PictureGenerator_l78_1 + 12'h007);
  assign _zz_when_PictureGenerator_l81_1_2 = {2'd0, coordinate_x};
  assign _zz_when_PictureGenerator_l87_1_1 = {2'd0, coordinate_x};
  assign _zz_when_PictureGenerator_l87_1_2 = {2'd0, coordinate_y};
  assign _zz_when_PictureGenerator_l87_1_3 = {2'd0, coordinate_x};
  assign _zz_when_PictureGenerator_l87_1_4 = (_zz_when_PictureGenerator_l78_1 + 12'h018);
  assign _zz_when_PictureGenerator_l87_1_5 = {2'd0, coordinate_y};
  assign _zz_when_PictureGenerator_l87_1_6 = (_zz_when_PictureGenerator_l87_1 + 12'h018);
  assign _zz_when_PictureGenerator_l138_1_1 = _zz_when_PictureGenerator_l138_3[2:0];
  assign _zz__zz_when_PictureGenerator_l138_5_1 = (_zz__zz_when_PictureGenerator_l138_5_2 + _zz_when_PictureGenerator_l78_2);
  assign _zz__zz_when_PictureGenerator_l138_5_3 = (10'h007 - coordinate_x);
  assign _zz__zz_when_PictureGenerator_l138_5_2 = {2'd0, _zz__zz_when_PictureGenerator_l138_5_3};
  assign _zz__zz_when_PictureGenerator_l138_4_3 = (_zz__zz_when_PictureGenerator_l138_4_4 - _zz_when_PictureGenerator_l87_2);
  assign _zz__zz_when_PictureGenerator_l138_4_2 = _zz__zz_when_PictureGenerator_l138_4_3[6:0];
  assign _zz__zz_when_PictureGenerator_l138_4_4 = (_zz__zz_when_PictureGenerator_l138_4_5 - _zz_when_PictureGenerator_l87_2);
  assign _zz__zz_when_PictureGenerator_l138_4_5 = (_zz__zz_when_PictureGenerator_l138_4_6 - _zz_when_PictureGenerator_l87_2);
  assign _zz__zz_when_PictureGenerator_l138_4_7 = (_zz__zz_when_PictureGenerator_l138_4_8 + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_4_6 = {2'd0, _zz__zz_when_PictureGenerator_l138_4_7};
  assign _zz__zz_when_PictureGenerator_l138_4_8 = (coordinate_y + coordinate_y);
  assign _zz_when_PictureGenerator_l78_2_1 = (_zz_when_PictureGenerator_l78_2 + 12'h00f);
  assign _zz_when_PictureGenerator_l78_2_2 = {2'd0, coordinate_x};
  assign _zz__zz_when_PictureGenerator_l138_5_4 = (_zz__zz_when_PictureGenerator_l138_5_5 + _zz_when_PictureGenerator_l78_2);
  assign _zz__zz_when_PictureGenerator_l138_5_6 = (10'h017 - coordinate_x);
  assign _zz__zz_when_PictureGenerator_l138_5_5 = {2'd0, _zz__zz_when_PictureGenerator_l138_5_6};
  assign _zz__zz_when_PictureGenerator_l138_4_11 = (12'h002 + _zz__zz_when_PictureGenerator_l138_4_12);
  assign _zz__zz_when_PictureGenerator_l138_4_10 = _zz__zz_when_PictureGenerator_l138_4_11[6:0];
  assign _zz__zz_when_PictureGenerator_l138_4_12 = (_zz__zz_when_PictureGenerator_l138_4_13 - _zz_when_PictureGenerator_l87_2);
  assign _zz__zz_when_PictureGenerator_l138_4_13 = (_zz__zz_when_PictureGenerator_l138_4_14 - _zz_when_PictureGenerator_l87_2);
  assign _zz__zz_when_PictureGenerator_l138_4_14 = (_zz__zz_when_PictureGenerator_l138_4_15 - _zz_when_PictureGenerator_l87_2);
  assign _zz__zz_when_PictureGenerator_l138_4_16 = (_zz__zz_when_PictureGenerator_l138_4_17 + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_4_15 = {2'd0, _zz__zz_when_PictureGenerator_l138_4_16};
  assign _zz__zz_when_PictureGenerator_l138_4_17 = (coordinate_y + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_5_7 = (_zz__zz_when_PictureGenerator_l138_5_8 + _zz_when_PictureGenerator_l78_2);
  assign _zz__zz_when_PictureGenerator_l138_5_9 = (10'h00f - coordinate_x);
  assign _zz__zz_when_PictureGenerator_l138_5_8 = {2'd0, _zz__zz_when_PictureGenerator_l138_5_9};
  assign _zz__zz_when_PictureGenerator_l138_4_20 = (12'h001 + _zz__zz_when_PictureGenerator_l138_4_21);
  assign _zz__zz_when_PictureGenerator_l138_4_19 = _zz__zz_when_PictureGenerator_l138_4_20[6:0];
  assign _zz__zz_when_PictureGenerator_l138_4_21 = (_zz__zz_when_PictureGenerator_l138_4_22 - _zz_when_PictureGenerator_l87_2);
  assign _zz__zz_when_PictureGenerator_l138_4_22 = (_zz__zz_when_PictureGenerator_l138_4_23 - _zz_when_PictureGenerator_l87_2);
  assign _zz__zz_when_PictureGenerator_l138_4_23 = (_zz__zz_when_PictureGenerator_l138_4_24 - _zz_when_PictureGenerator_l87_2);
  assign _zz__zz_when_PictureGenerator_l138_4_25 = (_zz__zz_when_PictureGenerator_l138_4_26 + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_4_24 = {2'd0, _zz__zz_when_PictureGenerator_l138_4_25};
  assign _zz__zz_when_PictureGenerator_l138_4_26 = (coordinate_y + coordinate_y);
  assign _zz_when_PictureGenerator_l81_2 = (_zz_when_PictureGenerator_l78_2 + 12'h007);
  assign _zz_when_PictureGenerator_l81_2_1 = {2'd0, coordinate_x};
  assign _zz_when_PictureGenerator_l87_2_1 = {2'd0, coordinate_x};
  assign _zz_when_PictureGenerator_l87_2_2 = {2'd0, coordinate_y};
  assign _zz_when_PictureGenerator_l87_2_3 = {2'd0, coordinate_x};
  assign _zz_when_PictureGenerator_l87_2_4 = (_zz_when_PictureGenerator_l78_2 + 12'h018);
  assign _zz_when_PictureGenerator_l87_2_5 = {2'd0, coordinate_y};
  assign _zz_when_PictureGenerator_l87_2_6 = (_zz_when_PictureGenerator_l87_2 + 12'h018);
  assign _zz_when_PictureGenerator_l138_2_1 = _zz_when_PictureGenerator_l138_5[2:0];
  assign _zz__zz_when_PictureGenerator_l138_7_1 = (_zz__zz_when_PictureGenerator_l138_7_2 + _zz_when_PictureGenerator_l78_3);
  assign _zz__zz_when_PictureGenerator_l138_7_3 = (10'h007 - coordinate_x);
  assign _zz__zz_when_PictureGenerator_l138_7_2 = {2'd0, _zz__zz_when_PictureGenerator_l138_7_3};
  assign _zz__zz_when_PictureGenerator_l138_6_3 = (_zz__zz_when_PictureGenerator_l138_6_4 - _zz_when_PictureGenerator_l87_3);
  assign _zz__zz_when_PictureGenerator_l138_6_2 = _zz__zz_when_PictureGenerator_l138_6_3[6:0];
  assign _zz__zz_when_PictureGenerator_l138_6_4 = (_zz__zz_when_PictureGenerator_l138_6_5 - _zz_when_PictureGenerator_l87_3);
  assign _zz__zz_when_PictureGenerator_l138_6_5 = (_zz__zz_when_PictureGenerator_l138_6_6 - _zz_when_PictureGenerator_l87_3);
  assign _zz__zz_when_PictureGenerator_l138_6_7 = (_zz__zz_when_PictureGenerator_l138_6_8 + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_6_6 = {2'd0, _zz__zz_when_PictureGenerator_l138_6_7};
  assign _zz__zz_when_PictureGenerator_l138_6_8 = (coordinate_y + coordinate_y);
  assign _zz_when_PictureGenerator_l78_3_1 = (_zz_when_PictureGenerator_l78_3 + 12'h00f);
  assign _zz_when_PictureGenerator_l78_3_2 = {2'd0, coordinate_x};
  assign _zz__zz_when_PictureGenerator_l138_7_4 = (_zz__zz_when_PictureGenerator_l138_7_5 + _zz_when_PictureGenerator_l78_3);
  assign _zz__zz_when_PictureGenerator_l138_7_6 = (10'h017 - coordinate_x);
  assign _zz__zz_when_PictureGenerator_l138_7_5 = {2'd0, _zz__zz_when_PictureGenerator_l138_7_6};
  assign _zz__zz_when_PictureGenerator_l138_6_11 = (12'h002 + _zz__zz_when_PictureGenerator_l138_6_12);
  assign _zz__zz_when_PictureGenerator_l138_6_10 = _zz__zz_when_PictureGenerator_l138_6_11[6:0];
  assign _zz__zz_when_PictureGenerator_l138_6_12 = (_zz__zz_when_PictureGenerator_l138_6_13 - _zz_when_PictureGenerator_l87_3);
  assign _zz__zz_when_PictureGenerator_l138_6_13 = (_zz__zz_when_PictureGenerator_l138_6_14 - _zz_when_PictureGenerator_l87_3);
  assign _zz__zz_when_PictureGenerator_l138_6_14 = (_zz__zz_when_PictureGenerator_l138_6_15 - _zz_when_PictureGenerator_l87_3);
  assign _zz__zz_when_PictureGenerator_l138_6_16 = (_zz__zz_when_PictureGenerator_l138_6_17 + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_6_15 = {2'd0, _zz__zz_when_PictureGenerator_l138_6_16};
  assign _zz__zz_when_PictureGenerator_l138_6_17 = (coordinate_y + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_7_7 = (_zz__zz_when_PictureGenerator_l138_7_8 + _zz_when_PictureGenerator_l78_3);
  assign _zz__zz_when_PictureGenerator_l138_7_9 = (10'h00f - coordinate_x);
  assign _zz__zz_when_PictureGenerator_l138_7_8 = {2'd0, _zz__zz_when_PictureGenerator_l138_7_9};
  assign _zz__zz_when_PictureGenerator_l138_6_20 = (12'h001 + _zz__zz_when_PictureGenerator_l138_6_21);
  assign _zz__zz_when_PictureGenerator_l138_6_19 = _zz__zz_when_PictureGenerator_l138_6_20[6:0];
  assign _zz__zz_when_PictureGenerator_l138_6_21 = (_zz__zz_when_PictureGenerator_l138_6_22 - _zz_when_PictureGenerator_l87_3);
  assign _zz__zz_when_PictureGenerator_l138_6_22 = (_zz__zz_when_PictureGenerator_l138_6_23 - _zz_when_PictureGenerator_l87_3);
  assign _zz__zz_when_PictureGenerator_l138_6_23 = (_zz__zz_when_PictureGenerator_l138_6_24 - _zz_when_PictureGenerator_l87_3);
  assign _zz__zz_when_PictureGenerator_l138_6_25 = (_zz__zz_when_PictureGenerator_l138_6_26 + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_6_24 = {2'd0, _zz__zz_when_PictureGenerator_l138_6_25};
  assign _zz__zz_when_PictureGenerator_l138_6_26 = (coordinate_y + coordinate_y);
  assign _zz_when_PictureGenerator_l81_3 = (_zz_when_PictureGenerator_l78_3 + 12'h007);
  assign _zz_when_PictureGenerator_l81_3_1 = {2'd0, coordinate_x};
  assign _zz_when_PictureGenerator_l87_3_1 = {2'd0, coordinate_x};
  assign _zz_when_PictureGenerator_l87_3_2 = {2'd0, coordinate_y};
  assign _zz_when_PictureGenerator_l87_3_3 = {2'd0, coordinate_x};
  assign _zz_when_PictureGenerator_l87_3_4 = (_zz_when_PictureGenerator_l78_3 + 12'h018);
  assign _zz_when_PictureGenerator_l87_3_5 = {2'd0, coordinate_y};
  assign _zz_when_PictureGenerator_l87_3_6 = (_zz_when_PictureGenerator_l87_3 + 12'h018);
  assign _zz_when_PictureGenerator_l138_3_1 = _zz_when_PictureGenerator_l138_7[2:0];
  assign _zz__zz_when_PictureGenerator_l138_9_1 = (_zz__zz_when_PictureGenerator_l138_9_2 + _zz_when_PictureGenerator_l78_4);
  assign _zz__zz_when_PictureGenerator_l138_9_3 = (10'h007 - coordinate_x);
  assign _zz__zz_when_PictureGenerator_l138_9_2 = {2'd0, _zz__zz_when_PictureGenerator_l138_9_3};
  assign _zz__zz_when_PictureGenerator_l138_8_3 = (_zz__zz_when_PictureGenerator_l138_8_4 - _zz_when_PictureGenerator_l87_4);
  assign _zz__zz_when_PictureGenerator_l138_8_2 = _zz__zz_when_PictureGenerator_l138_8_3[6:0];
  assign _zz__zz_when_PictureGenerator_l138_8_4 = (_zz__zz_when_PictureGenerator_l138_8_5 - _zz_when_PictureGenerator_l87_4);
  assign _zz__zz_when_PictureGenerator_l138_8_5 = (_zz__zz_when_PictureGenerator_l138_8_6 - _zz_when_PictureGenerator_l87_4);
  assign _zz__zz_when_PictureGenerator_l138_8_7 = (_zz__zz_when_PictureGenerator_l138_8_8 + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_8_6 = {2'd0, _zz__zz_when_PictureGenerator_l138_8_7};
  assign _zz__zz_when_PictureGenerator_l138_8_8 = (coordinate_y + coordinate_y);
  assign _zz_when_PictureGenerator_l78_4_1 = (_zz_when_PictureGenerator_l78_4 + 12'h00f);
  assign _zz_when_PictureGenerator_l78_4_2 = {2'd0, coordinate_x};
  assign _zz__zz_when_PictureGenerator_l138_9_4 = (_zz__zz_when_PictureGenerator_l138_9_5 + _zz_when_PictureGenerator_l78_4);
  assign _zz__zz_when_PictureGenerator_l138_9_6 = (10'h017 - coordinate_x);
  assign _zz__zz_when_PictureGenerator_l138_9_5 = {2'd0, _zz__zz_when_PictureGenerator_l138_9_6};
  assign _zz__zz_when_PictureGenerator_l138_8_11 = (12'h002 + _zz__zz_when_PictureGenerator_l138_8_12);
  assign _zz__zz_when_PictureGenerator_l138_8_10 = _zz__zz_when_PictureGenerator_l138_8_11[6:0];
  assign _zz__zz_when_PictureGenerator_l138_8_12 = (_zz__zz_when_PictureGenerator_l138_8_13 - _zz_when_PictureGenerator_l87_4);
  assign _zz__zz_when_PictureGenerator_l138_8_13 = (_zz__zz_when_PictureGenerator_l138_8_14 - _zz_when_PictureGenerator_l87_4);
  assign _zz__zz_when_PictureGenerator_l138_8_14 = (_zz__zz_when_PictureGenerator_l138_8_15 - _zz_when_PictureGenerator_l87_4);
  assign _zz__zz_when_PictureGenerator_l138_8_16 = (_zz__zz_when_PictureGenerator_l138_8_17 + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_8_15 = {2'd0, _zz__zz_when_PictureGenerator_l138_8_16};
  assign _zz__zz_when_PictureGenerator_l138_8_17 = (coordinate_y + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_9_7 = (_zz__zz_when_PictureGenerator_l138_9_8 + _zz_when_PictureGenerator_l78_4);
  assign _zz__zz_when_PictureGenerator_l138_9_9 = (10'h00f - coordinate_x);
  assign _zz__zz_when_PictureGenerator_l138_9_8 = {2'd0, _zz__zz_when_PictureGenerator_l138_9_9};
  assign _zz__zz_when_PictureGenerator_l138_8_20 = (12'h001 + _zz__zz_when_PictureGenerator_l138_8_21);
  assign _zz__zz_when_PictureGenerator_l138_8_19 = _zz__zz_when_PictureGenerator_l138_8_20[6:0];
  assign _zz__zz_when_PictureGenerator_l138_8_21 = (_zz__zz_when_PictureGenerator_l138_8_22 - _zz_when_PictureGenerator_l87_4);
  assign _zz__zz_when_PictureGenerator_l138_8_22 = (_zz__zz_when_PictureGenerator_l138_8_23 - _zz_when_PictureGenerator_l87_4);
  assign _zz__zz_when_PictureGenerator_l138_8_23 = (_zz__zz_when_PictureGenerator_l138_8_24 - _zz_when_PictureGenerator_l87_4);
  assign _zz__zz_when_PictureGenerator_l138_8_25 = (_zz__zz_when_PictureGenerator_l138_8_26 + coordinate_y);
  assign _zz__zz_when_PictureGenerator_l138_8_24 = {2'd0, _zz__zz_when_PictureGenerator_l138_8_25};
  assign _zz__zz_when_PictureGenerator_l138_8_26 = (coordinate_y + coordinate_y);
  assign _zz_when_PictureGenerator_l81_4 = (_zz_when_PictureGenerator_l78_4 + 12'h007);
  assign _zz_when_PictureGenerator_l81_4_1 = {2'd0, coordinate_x};
  assign _zz_when_PictureGenerator_l87_4_1 = {2'd0, coordinate_x};
  assign _zz_when_PictureGenerator_l87_4_2 = {2'd0, coordinate_y};
  assign _zz_when_PictureGenerator_l87_4_3 = {2'd0, coordinate_x};
  assign _zz_when_PictureGenerator_l87_4_4 = (_zz_when_PictureGenerator_l78_4 + 12'h018);
  assign _zz_when_PictureGenerator_l87_4_5 = {2'd0, coordinate_y};
  assign _zz_when_PictureGenerator_l87_4_6 = (_zz_when_PictureGenerator_l87_4 + 12'h018);
  assign _zz_when_PictureGenerator_l138_4_1 = _zz_when_PictureGenerator_l138_9[2:0];
  RAddressGen rAddr (
    .ram_en   (rAddr_ram_en[4:0]   ), //o
    .ram_x    (rAddr_ram_x[9:0]    ), //i
    .ram_y    (rAddr_ram_y[9:0]    ), //i
    .ram_addr (rAddr_ram_addr[13:0]), //o
    .clk      (clk                 ), //i
    .reset    (reset               )  //i
  );
  always @(*) begin
    case(_zz__zz_when_PictureGenerator_l138_2)
      7'b0000000 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_0;
      7'b0000001 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_1;
      7'b0000010 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_2;
      7'b0000011 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_3;
      7'b0000100 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_4;
      7'b0000101 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_5;
      7'b0000110 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_6;
      7'b0000111 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_7;
      7'b0001000 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_8;
      7'b0001001 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_9;
      7'b0001010 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_10;
      7'b0001011 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_11;
      7'b0001100 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_12;
      7'b0001101 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_13;
      7'b0001110 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_14;
      7'b0001111 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_15;
      7'b0010000 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_16;
      7'b0010001 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_17;
      7'b0010010 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_18;
      7'b0010011 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_19;
      7'b0010100 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_20;
      7'b0010101 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_21;
      7'b0010110 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_22;
      7'b0010111 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_23;
      7'b0011000 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_24;
      7'b0011001 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_25;
      7'b0011010 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_26;
      7'b0011011 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_27;
      7'b0011100 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_28;
      7'b0011101 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_29;
      7'b0011110 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_30;
      7'b0011111 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_31;
      7'b0100000 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_32;
      7'b0100001 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_33;
      7'b0100010 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_34;
      7'b0100011 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_35;
      7'b0100100 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_36;
      7'b0100101 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_37;
      7'b0100110 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_38;
      7'b0100111 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_39;
      7'b0101000 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_40;
      7'b0101001 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_41;
      7'b0101010 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_42;
      7'b0101011 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_43;
      7'b0101100 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_44;
      7'b0101101 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_45;
      7'b0101110 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_46;
      7'b0101111 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_47;
      7'b0110000 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_48;
      7'b0110001 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_49;
      7'b0110010 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_50;
      7'b0110011 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_51;
      7'b0110100 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_52;
      7'b0110101 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_53;
      7'b0110110 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_54;
      7'b0110111 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_55;
      7'b0111000 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_56;
      7'b0111001 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_57;
      7'b0111010 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_58;
      7'b0111011 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_59;
      7'b0111100 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_60;
      7'b0111101 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_61;
      7'b0111110 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_62;
      7'b0111111 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_63;
      7'b1000000 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_64;
      7'b1000001 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_65;
      7'b1000010 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_66;
      7'b1000011 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_67;
      7'b1000100 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_68;
      7'b1000101 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_69;
      7'b1000110 : _zz__zz_when_PictureGenerator_l138 = fontVec_0_70;
      default : _zz__zz_when_PictureGenerator_l138 = fontVec_0_71;
    endcase
  end

  always @(*) begin
    case(_zz__zz_when_PictureGenerator_l138_10)
      7'b0000000 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_0;
      7'b0000001 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_1;
      7'b0000010 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_2;
      7'b0000011 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_3;
      7'b0000100 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_4;
      7'b0000101 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_5;
      7'b0000110 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_6;
      7'b0000111 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_7;
      7'b0001000 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_8;
      7'b0001001 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_9;
      7'b0001010 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_10;
      7'b0001011 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_11;
      7'b0001100 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_12;
      7'b0001101 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_13;
      7'b0001110 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_14;
      7'b0001111 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_15;
      7'b0010000 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_16;
      7'b0010001 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_17;
      7'b0010010 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_18;
      7'b0010011 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_19;
      7'b0010100 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_20;
      7'b0010101 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_21;
      7'b0010110 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_22;
      7'b0010111 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_23;
      7'b0011000 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_24;
      7'b0011001 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_25;
      7'b0011010 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_26;
      7'b0011011 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_27;
      7'b0011100 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_28;
      7'b0011101 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_29;
      7'b0011110 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_30;
      7'b0011111 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_31;
      7'b0100000 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_32;
      7'b0100001 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_33;
      7'b0100010 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_34;
      7'b0100011 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_35;
      7'b0100100 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_36;
      7'b0100101 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_37;
      7'b0100110 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_38;
      7'b0100111 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_39;
      7'b0101000 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_40;
      7'b0101001 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_41;
      7'b0101010 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_42;
      7'b0101011 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_43;
      7'b0101100 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_44;
      7'b0101101 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_45;
      7'b0101110 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_46;
      7'b0101111 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_47;
      7'b0110000 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_48;
      7'b0110001 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_49;
      7'b0110010 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_50;
      7'b0110011 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_51;
      7'b0110100 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_52;
      7'b0110101 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_53;
      7'b0110110 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_54;
      7'b0110111 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_55;
      7'b0111000 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_56;
      7'b0111001 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_57;
      7'b0111010 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_58;
      7'b0111011 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_59;
      7'b0111100 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_60;
      7'b0111101 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_61;
      7'b0111110 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_62;
      7'b0111111 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_63;
      7'b1000000 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_64;
      7'b1000001 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_65;
      7'b1000010 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_66;
      7'b1000011 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_67;
      7'b1000100 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_68;
      7'b1000101 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_69;
      7'b1000110 : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_70;
      default : _zz__zz_when_PictureGenerator_l138_9 = fontVec_0_71;
    endcase
  end

  always @(*) begin
    case(_zz__zz_when_PictureGenerator_l138_19)
      7'b0000000 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_0;
      7'b0000001 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_1;
      7'b0000010 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_2;
      7'b0000011 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_3;
      7'b0000100 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_4;
      7'b0000101 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_5;
      7'b0000110 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_6;
      7'b0000111 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_7;
      7'b0001000 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_8;
      7'b0001001 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_9;
      7'b0001010 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_10;
      7'b0001011 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_11;
      7'b0001100 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_12;
      7'b0001101 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_13;
      7'b0001110 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_14;
      7'b0001111 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_15;
      7'b0010000 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_16;
      7'b0010001 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_17;
      7'b0010010 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_18;
      7'b0010011 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_19;
      7'b0010100 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_20;
      7'b0010101 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_21;
      7'b0010110 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_22;
      7'b0010111 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_23;
      7'b0011000 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_24;
      7'b0011001 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_25;
      7'b0011010 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_26;
      7'b0011011 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_27;
      7'b0011100 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_28;
      7'b0011101 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_29;
      7'b0011110 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_30;
      7'b0011111 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_31;
      7'b0100000 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_32;
      7'b0100001 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_33;
      7'b0100010 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_34;
      7'b0100011 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_35;
      7'b0100100 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_36;
      7'b0100101 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_37;
      7'b0100110 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_38;
      7'b0100111 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_39;
      7'b0101000 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_40;
      7'b0101001 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_41;
      7'b0101010 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_42;
      7'b0101011 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_43;
      7'b0101100 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_44;
      7'b0101101 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_45;
      7'b0101110 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_46;
      7'b0101111 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_47;
      7'b0110000 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_48;
      7'b0110001 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_49;
      7'b0110010 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_50;
      7'b0110011 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_51;
      7'b0110100 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_52;
      7'b0110101 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_53;
      7'b0110110 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_54;
      7'b0110111 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_55;
      7'b0111000 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_56;
      7'b0111001 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_57;
      7'b0111010 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_58;
      7'b0111011 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_59;
      7'b0111100 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_60;
      7'b0111101 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_61;
      7'b0111110 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_62;
      7'b0111111 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_63;
      7'b1000000 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_64;
      7'b1000001 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_65;
      7'b1000010 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_66;
      7'b1000011 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_67;
      7'b1000100 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_68;
      7'b1000101 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_69;
      7'b1000110 : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_70;
      default : _zz__zz_when_PictureGenerator_l138_18 = fontVec_0_71;
    endcase
  end

  always @(*) begin
    case(_zz__zz_when_PictureGenerator_l138_2_2)
      7'b0000000 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_0;
      7'b0000001 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_1;
      7'b0000010 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_2;
      7'b0000011 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_3;
      7'b0000100 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_4;
      7'b0000101 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_5;
      7'b0000110 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_6;
      7'b0000111 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_7;
      7'b0001000 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_8;
      7'b0001001 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_9;
      7'b0001010 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_10;
      7'b0001011 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_11;
      7'b0001100 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_12;
      7'b0001101 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_13;
      7'b0001110 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_14;
      7'b0001111 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_15;
      7'b0010000 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_16;
      7'b0010001 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_17;
      7'b0010010 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_18;
      7'b0010011 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_19;
      7'b0010100 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_20;
      7'b0010101 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_21;
      7'b0010110 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_22;
      7'b0010111 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_23;
      7'b0011000 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_24;
      7'b0011001 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_25;
      7'b0011010 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_26;
      7'b0011011 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_27;
      7'b0011100 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_28;
      7'b0011101 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_29;
      7'b0011110 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_30;
      7'b0011111 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_31;
      7'b0100000 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_32;
      7'b0100001 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_33;
      7'b0100010 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_34;
      7'b0100011 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_35;
      7'b0100100 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_36;
      7'b0100101 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_37;
      7'b0100110 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_38;
      7'b0100111 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_39;
      7'b0101000 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_40;
      7'b0101001 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_41;
      7'b0101010 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_42;
      7'b0101011 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_43;
      7'b0101100 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_44;
      7'b0101101 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_45;
      7'b0101110 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_46;
      7'b0101111 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_47;
      7'b0110000 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_48;
      7'b0110001 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_49;
      7'b0110010 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_50;
      7'b0110011 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_51;
      7'b0110100 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_52;
      7'b0110101 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_53;
      7'b0110110 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_54;
      7'b0110111 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_55;
      7'b0111000 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_56;
      7'b0111001 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_57;
      7'b0111010 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_58;
      7'b0111011 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_59;
      7'b0111100 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_60;
      7'b0111101 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_61;
      7'b0111110 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_62;
      7'b0111111 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_63;
      7'b1000000 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_64;
      7'b1000001 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_65;
      7'b1000010 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_66;
      7'b1000011 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_67;
      7'b1000100 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_68;
      7'b1000101 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_69;
      7'b1000110 : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_70;
      default : _zz__zz_when_PictureGenerator_l138_2_1 = fontVec_1_71;
    endcase
  end

  always @(*) begin
    case(_zz__zz_when_PictureGenerator_l138_2_10)
      7'b0000000 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_0;
      7'b0000001 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_1;
      7'b0000010 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_2;
      7'b0000011 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_3;
      7'b0000100 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_4;
      7'b0000101 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_5;
      7'b0000110 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_6;
      7'b0000111 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_7;
      7'b0001000 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_8;
      7'b0001001 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_9;
      7'b0001010 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_10;
      7'b0001011 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_11;
      7'b0001100 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_12;
      7'b0001101 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_13;
      7'b0001110 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_14;
      7'b0001111 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_15;
      7'b0010000 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_16;
      7'b0010001 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_17;
      7'b0010010 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_18;
      7'b0010011 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_19;
      7'b0010100 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_20;
      7'b0010101 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_21;
      7'b0010110 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_22;
      7'b0010111 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_23;
      7'b0011000 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_24;
      7'b0011001 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_25;
      7'b0011010 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_26;
      7'b0011011 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_27;
      7'b0011100 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_28;
      7'b0011101 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_29;
      7'b0011110 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_30;
      7'b0011111 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_31;
      7'b0100000 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_32;
      7'b0100001 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_33;
      7'b0100010 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_34;
      7'b0100011 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_35;
      7'b0100100 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_36;
      7'b0100101 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_37;
      7'b0100110 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_38;
      7'b0100111 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_39;
      7'b0101000 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_40;
      7'b0101001 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_41;
      7'b0101010 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_42;
      7'b0101011 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_43;
      7'b0101100 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_44;
      7'b0101101 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_45;
      7'b0101110 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_46;
      7'b0101111 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_47;
      7'b0110000 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_48;
      7'b0110001 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_49;
      7'b0110010 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_50;
      7'b0110011 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_51;
      7'b0110100 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_52;
      7'b0110101 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_53;
      7'b0110110 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_54;
      7'b0110111 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_55;
      7'b0111000 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_56;
      7'b0111001 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_57;
      7'b0111010 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_58;
      7'b0111011 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_59;
      7'b0111100 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_60;
      7'b0111101 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_61;
      7'b0111110 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_62;
      7'b0111111 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_63;
      7'b1000000 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_64;
      7'b1000001 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_65;
      7'b1000010 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_66;
      7'b1000011 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_67;
      7'b1000100 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_68;
      7'b1000101 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_69;
      7'b1000110 : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_70;
      default : _zz__zz_when_PictureGenerator_l138_2_9 = fontVec_1_71;
    endcase
  end

  always @(*) begin
    case(_zz__zz_when_PictureGenerator_l138_2_19)
      7'b0000000 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_0;
      7'b0000001 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_1;
      7'b0000010 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_2;
      7'b0000011 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_3;
      7'b0000100 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_4;
      7'b0000101 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_5;
      7'b0000110 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_6;
      7'b0000111 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_7;
      7'b0001000 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_8;
      7'b0001001 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_9;
      7'b0001010 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_10;
      7'b0001011 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_11;
      7'b0001100 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_12;
      7'b0001101 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_13;
      7'b0001110 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_14;
      7'b0001111 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_15;
      7'b0010000 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_16;
      7'b0010001 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_17;
      7'b0010010 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_18;
      7'b0010011 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_19;
      7'b0010100 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_20;
      7'b0010101 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_21;
      7'b0010110 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_22;
      7'b0010111 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_23;
      7'b0011000 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_24;
      7'b0011001 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_25;
      7'b0011010 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_26;
      7'b0011011 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_27;
      7'b0011100 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_28;
      7'b0011101 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_29;
      7'b0011110 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_30;
      7'b0011111 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_31;
      7'b0100000 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_32;
      7'b0100001 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_33;
      7'b0100010 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_34;
      7'b0100011 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_35;
      7'b0100100 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_36;
      7'b0100101 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_37;
      7'b0100110 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_38;
      7'b0100111 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_39;
      7'b0101000 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_40;
      7'b0101001 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_41;
      7'b0101010 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_42;
      7'b0101011 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_43;
      7'b0101100 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_44;
      7'b0101101 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_45;
      7'b0101110 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_46;
      7'b0101111 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_47;
      7'b0110000 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_48;
      7'b0110001 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_49;
      7'b0110010 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_50;
      7'b0110011 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_51;
      7'b0110100 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_52;
      7'b0110101 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_53;
      7'b0110110 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_54;
      7'b0110111 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_55;
      7'b0111000 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_56;
      7'b0111001 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_57;
      7'b0111010 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_58;
      7'b0111011 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_59;
      7'b0111100 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_60;
      7'b0111101 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_61;
      7'b0111110 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_62;
      7'b0111111 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_63;
      7'b1000000 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_64;
      7'b1000001 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_65;
      7'b1000010 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_66;
      7'b1000011 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_67;
      7'b1000100 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_68;
      7'b1000101 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_69;
      7'b1000110 : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_70;
      default : _zz__zz_when_PictureGenerator_l138_2_18 = fontVec_1_71;
    endcase
  end

  always @(*) begin
    case(_zz__zz_when_PictureGenerator_l138_4_2)
      7'b0000000 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_0;
      7'b0000001 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_1;
      7'b0000010 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_2;
      7'b0000011 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_3;
      7'b0000100 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_4;
      7'b0000101 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_5;
      7'b0000110 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_6;
      7'b0000111 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_7;
      7'b0001000 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_8;
      7'b0001001 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_9;
      7'b0001010 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_10;
      7'b0001011 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_11;
      7'b0001100 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_12;
      7'b0001101 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_13;
      7'b0001110 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_14;
      7'b0001111 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_15;
      7'b0010000 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_16;
      7'b0010001 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_17;
      7'b0010010 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_18;
      7'b0010011 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_19;
      7'b0010100 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_20;
      7'b0010101 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_21;
      7'b0010110 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_22;
      7'b0010111 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_23;
      7'b0011000 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_24;
      7'b0011001 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_25;
      7'b0011010 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_26;
      7'b0011011 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_27;
      7'b0011100 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_28;
      7'b0011101 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_29;
      7'b0011110 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_30;
      7'b0011111 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_31;
      7'b0100000 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_32;
      7'b0100001 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_33;
      7'b0100010 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_34;
      7'b0100011 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_35;
      7'b0100100 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_36;
      7'b0100101 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_37;
      7'b0100110 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_38;
      7'b0100111 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_39;
      7'b0101000 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_40;
      7'b0101001 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_41;
      7'b0101010 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_42;
      7'b0101011 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_43;
      7'b0101100 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_44;
      7'b0101101 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_45;
      7'b0101110 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_46;
      7'b0101111 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_47;
      7'b0110000 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_48;
      7'b0110001 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_49;
      7'b0110010 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_50;
      7'b0110011 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_51;
      7'b0110100 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_52;
      7'b0110101 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_53;
      7'b0110110 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_54;
      7'b0110111 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_55;
      7'b0111000 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_56;
      7'b0111001 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_57;
      7'b0111010 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_58;
      7'b0111011 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_59;
      7'b0111100 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_60;
      7'b0111101 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_61;
      7'b0111110 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_62;
      7'b0111111 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_63;
      7'b1000000 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_64;
      7'b1000001 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_65;
      7'b1000010 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_66;
      7'b1000011 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_67;
      7'b1000100 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_68;
      7'b1000101 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_69;
      7'b1000110 : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_70;
      default : _zz__zz_when_PictureGenerator_l138_4_1 = fontVec_2_71;
    endcase
  end

  always @(*) begin
    case(_zz__zz_when_PictureGenerator_l138_4_10)
      7'b0000000 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_0;
      7'b0000001 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_1;
      7'b0000010 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_2;
      7'b0000011 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_3;
      7'b0000100 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_4;
      7'b0000101 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_5;
      7'b0000110 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_6;
      7'b0000111 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_7;
      7'b0001000 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_8;
      7'b0001001 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_9;
      7'b0001010 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_10;
      7'b0001011 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_11;
      7'b0001100 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_12;
      7'b0001101 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_13;
      7'b0001110 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_14;
      7'b0001111 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_15;
      7'b0010000 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_16;
      7'b0010001 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_17;
      7'b0010010 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_18;
      7'b0010011 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_19;
      7'b0010100 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_20;
      7'b0010101 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_21;
      7'b0010110 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_22;
      7'b0010111 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_23;
      7'b0011000 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_24;
      7'b0011001 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_25;
      7'b0011010 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_26;
      7'b0011011 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_27;
      7'b0011100 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_28;
      7'b0011101 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_29;
      7'b0011110 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_30;
      7'b0011111 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_31;
      7'b0100000 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_32;
      7'b0100001 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_33;
      7'b0100010 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_34;
      7'b0100011 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_35;
      7'b0100100 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_36;
      7'b0100101 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_37;
      7'b0100110 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_38;
      7'b0100111 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_39;
      7'b0101000 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_40;
      7'b0101001 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_41;
      7'b0101010 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_42;
      7'b0101011 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_43;
      7'b0101100 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_44;
      7'b0101101 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_45;
      7'b0101110 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_46;
      7'b0101111 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_47;
      7'b0110000 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_48;
      7'b0110001 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_49;
      7'b0110010 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_50;
      7'b0110011 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_51;
      7'b0110100 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_52;
      7'b0110101 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_53;
      7'b0110110 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_54;
      7'b0110111 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_55;
      7'b0111000 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_56;
      7'b0111001 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_57;
      7'b0111010 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_58;
      7'b0111011 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_59;
      7'b0111100 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_60;
      7'b0111101 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_61;
      7'b0111110 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_62;
      7'b0111111 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_63;
      7'b1000000 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_64;
      7'b1000001 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_65;
      7'b1000010 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_66;
      7'b1000011 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_67;
      7'b1000100 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_68;
      7'b1000101 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_69;
      7'b1000110 : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_70;
      default : _zz__zz_when_PictureGenerator_l138_4_9 = fontVec_2_71;
    endcase
  end

  always @(*) begin
    case(_zz__zz_when_PictureGenerator_l138_4_19)
      7'b0000000 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_0;
      7'b0000001 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_1;
      7'b0000010 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_2;
      7'b0000011 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_3;
      7'b0000100 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_4;
      7'b0000101 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_5;
      7'b0000110 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_6;
      7'b0000111 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_7;
      7'b0001000 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_8;
      7'b0001001 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_9;
      7'b0001010 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_10;
      7'b0001011 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_11;
      7'b0001100 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_12;
      7'b0001101 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_13;
      7'b0001110 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_14;
      7'b0001111 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_15;
      7'b0010000 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_16;
      7'b0010001 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_17;
      7'b0010010 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_18;
      7'b0010011 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_19;
      7'b0010100 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_20;
      7'b0010101 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_21;
      7'b0010110 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_22;
      7'b0010111 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_23;
      7'b0011000 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_24;
      7'b0011001 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_25;
      7'b0011010 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_26;
      7'b0011011 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_27;
      7'b0011100 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_28;
      7'b0011101 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_29;
      7'b0011110 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_30;
      7'b0011111 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_31;
      7'b0100000 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_32;
      7'b0100001 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_33;
      7'b0100010 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_34;
      7'b0100011 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_35;
      7'b0100100 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_36;
      7'b0100101 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_37;
      7'b0100110 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_38;
      7'b0100111 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_39;
      7'b0101000 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_40;
      7'b0101001 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_41;
      7'b0101010 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_42;
      7'b0101011 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_43;
      7'b0101100 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_44;
      7'b0101101 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_45;
      7'b0101110 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_46;
      7'b0101111 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_47;
      7'b0110000 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_48;
      7'b0110001 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_49;
      7'b0110010 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_50;
      7'b0110011 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_51;
      7'b0110100 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_52;
      7'b0110101 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_53;
      7'b0110110 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_54;
      7'b0110111 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_55;
      7'b0111000 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_56;
      7'b0111001 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_57;
      7'b0111010 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_58;
      7'b0111011 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_59;
      7'b0111100 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_60;
      7'b0111101 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_61;
      7'b0111110 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_62;
      7'b0111111 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_63;
      7'b1000000 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_64;
      7'b1000001 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_65;
      7'b1000010 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_66;
      7'b1000011 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_67;
      7'b1000100 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_68;
      7'b1000101 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_69;
      7'b1000110 : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_70;
      default : _zz__zz_when_PictureGenerator_l138_4_18 = fontVec_2_71;
    endcase
  end

  always @(*) begin
    case(_zz__zz_when_PictureGenerator_l138_6_2)
      7'b0000000 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_0;
      7'b0000001 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_1;
      7'b0000010 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_2;
      7'b0000011 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_3;
      7'b0000100 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_4;
      7'b0000101 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_5;
      7'b0000110 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_6;
      7'b0000111 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_7;
      7'b0001000 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_8;
      7'b0001001 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_9;
      7'b0001010 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_10;
      7'b0001011 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_11;
      7'b0001100 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_12;
      7'b0001101 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_13;
      7'b0001110 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_14;
      7'b0001111 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_15;
      7'b0010000 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_16;
      7'b0010001 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_17;
      7'b0010010 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_18;
      7'b0010011 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_19;
      7'b0010100 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_20;
      7'b0010101 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_21;
      7'b0010110 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_22;
      7'b0010111 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_23;
      7'b0011000 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_24;
      7'b0011001 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_25;
      7'b0011010 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_26;
      7'b0011011 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_27;
      7'b0011100 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_28;
      7'b0011101 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_29;
      7'b0011110 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_30;
      7'b0011111 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_31;
      7'b0100000 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_32;
      7'b0100001 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_33;
      7'b0100010 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_34;
      7'b0100011 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_35;
      7'b0100100 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_36;
      7'b0100101 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_37;
      7'b0100110 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_38;
      7'b0100111 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_39;
      7'b0101000 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_40;
      7'b0101001 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_41;
      7'b0101010 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_42;
      7'b0101011 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_43;
      7'b0101100 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_44;
      7'b0101101 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_45;
      7'b0101110 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_46;
      7'b0101111 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_47;
      7'b0110000 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_48;
      7'b0110001 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_49;
      7'b0110010 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_50;
      7'b0110011 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_51;
      7'b0110100 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_52;
      7'b0110101 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_53;
      7'b0110110 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_54;
      7'b0110111 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_55;
      7'b0111000 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_56;
      7'b0111001 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_57;
      7'b0111010 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_58;
      7'b0111011 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_59;
      7'b0111100 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_60;
      7'b0111101 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_61;
      7'b0111110 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_62;
      7'b0111111 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_63;
      7'b1000000 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_64;
      7'b1000001 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_65;
      7'b1000010 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_66;
      7'b1000011 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_67;
      7'b1000100 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_68;
      7'b1000101 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_69;
      7'b1000110 : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_70;
      default : _zz__zz_when_PictureGenerator_l138_6_1 = fontVec_3_71;
    endcase
  end

  always @(*) begin
    case(_zz__zz_when_PictureGenerator_l138_6_10)
      7'b0000000 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_0;
      7'b0000001 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_1;
      7'b0000010 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_2;
      7'b0000011 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_3;
      7'b0000100 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_4;
      7'b0000101 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_5;
      7'b0000110 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_6;
      7'b0000111 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_7;
      7'b0001000 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_8;
      7'b0001001 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_9;
      7'b0001010 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_10;
      7'b0001011 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_11;
      7'b0001100 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_12;
      7'b0001101 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_13;
      7'b0001110 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_14;
      7'b0001111 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_15;
      7'b0010000 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_16;
      7'b0010001 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_17;
      7'b0010010 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_18;
      7'b0010011 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_19;
      7'b0010100 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_20;
      7'b0010101 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_21;
      7'b0010110 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_22;
      7'b0010111 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_23;
      7'b0011000 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_24;
      7'b0011001 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_25;
      7'b0011010 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_26;
      7'b0011011 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_27;
      7'b0011100 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_28;
      7'b0011101 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_29;
      7'b0011110 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_30;
      7'b0011111 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_31;
      7'b0100000 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_32;
      7'b0100001 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_33;
      7'b0100010 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_34;
      7'b0100011 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_35;
      7'b0100100 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_36;
      7'b0100101 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_37;
      7'b0100110 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_38;
      7'b0100111 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_39;
      7'b0101000 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_40;
      7'b0101001 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_41;
      7'b0101010 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_42;
      7'b0101011 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_43;
      7'b0101100 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_44;
      7'b0101101 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_45;
      7'b0101110 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_46;
      7'b0101111 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_47;
      7'b0110000 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_48;
      7'b0110001 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_49;
      7'b0110010 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_50;
      7'b0110011 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_51;
      7'b0110100 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_52;
      7'b0110101 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_53;
      7'b0110110 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_54;
      7'b0110111 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_55;
      7'b0111000 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_56;
      7'b0111001 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_57;
      7'b0111010 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_58;
      7'b0111011 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_59;
      7'b0111100 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_60;
      7'b0111101 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_61;
      7'b0111110 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_62;
      7'b0111111 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_63;
      7'b1000000 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_64;
      7'b1000001 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_65;
      7'b1000010 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_66;
      7'b1000011 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_67;
      7'b1000100 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_68;
      7'b1000101 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_69;
      7'b1000110 : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_70;
      default : _zz__zz_when_PictureGenerator_l138_6_9 = fontVec_3_71;
    endcase
  end

  always @(*) begin
    case(_zz__zz_when_PictureGenerator_l138_6_19)
      7'b0000000 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_0;
      7'b0000001 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_1;
      7'b0000010 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_2;
      7'b0000011 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_3;
      7'b0000100 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_4;
      7'b0000101 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_5;
      7'b0000110 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_6;
      7'b0000111 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_7;
      7'b0001000 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_8;
      7'b0001001 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_9;
      7'b0001010 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_10;
      7'b0001011 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_11;
      7'b0001100 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_12;
      7'b0001101 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_13;
      7'b0001110 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_14;
      7'b0001111 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_15;
      7'b0010000 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_16;
      7'b0010001 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_17;
      7'b0010010 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_18;
      7'b0010011 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_19;
      7'b0010100 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_20;
      7'b0010101 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_21;
      7'b0010110 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_22;
      7'b0010111 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_23;
      7'b0011000 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_24;
      7'b0011001 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_25;
      7'b0011010 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_26;
      7'b0011011 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_27;
      7'b0011100 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_28;
      7'b0011101 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_29;
      7'b0011110 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_30;
      7'b0011111 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_31;
      7'b0100000 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_32;
      7'b0100001 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_33;
      7'b0100010 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_34;
      7'b0100011 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_35;
      7'b0100100 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_36;
      7'b0100101 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_37;
      7'b0100110 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_38;
      7'b0100111 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_39;
      7'b0101000 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_40;
      7'b0101001 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_41;
      7'b0101010 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_42;
      7'b0101011 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_43;
      7'b0101100 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_44;
      7'b0101101 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_45;
      7'b0101110 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_46;
      7'b0101111 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_47;
      7'b0110000 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_48;
      7'b0110001 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_49;
      7'b0110010 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_50;
      7'b0110011 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_51;
      7'b0110100 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_52;
      7'b0110101 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_53;
      7'b0110110 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_54;
      7'b0110111 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_55;
      7'b0111000 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_56;
      7'b0111001 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_57;
      7'b0111010 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_58;
      7'b0111011 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_59;
      7'b0111100 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_60;
      7'b0111101 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_61;
      7'b0111110 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_62;
      7'b0111111 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_63;
      7'b1000000 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_64;
      7'b1000001 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_65;
      7'b1000010 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_66;
      7'b1000011 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_67;
      7'b1000100 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_68;
      7'b1000101 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_69;
      7'b1000110 : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_70;
      default : _zz__zz_when_PictureGenerator_l138_6_18 = fontVec_3_71;
    endcase
  end

  always @(*) begin
    case(_zz__zz_when_PictureGenerator_l138_8_2)
      7'b0000000 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_0;
      7'b0000001 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_1;
      7'b0000010 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_2;
      7'b0000011 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_3;
      7'b0000100 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_4;
      7'b0000101 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_5;
      7'b0000110 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_6;
      7'b0000111 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_7;
      7'b0001000 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_8;
      7'b0001001 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_9;
      7'b0001010 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_10;
      7'b0001011 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_11;
      7'b0001100 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_12;
      7'b0001101 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_13;
      7'b0001110 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_14;
      7'b0001111 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_15;
      7'b0010000 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_16;
      7'b0010001 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_17;
      7'b0010010 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_18;
      7'b0010011 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_19;
      7'b0010100 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_20;
      7'b0010101 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_21;
      7'b0010110 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_22;
      7'b0010111 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_23;
      7'b0011000 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_24;
      7'b0011001 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_25;
      7'b0011010 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_26;
      7'b0011011 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_27;
      7'b0011100 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_28;
      7'b0011101 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_29;
      7'b0011110 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_30;
      7'b0011111 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_31;
      7'b0100000 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_32;
      7'b0100001 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_33;
      7'b0100010 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_34;
      7'b0100011 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_35;
      7'b0100100 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_36;
      7'b0100101 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_37;
      7'b0100110 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_38;
      7'b0100111 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_39;
      7'b0101000 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_40;
      7'b0101001 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_41;
      7'b0101010 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_42;
      7'b0101011 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_43;
      7'b0101100 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_44;
      7'b0101101 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_45;
      7'b0101110 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_46;
      7'b0101111 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_47;
      7'b0110000 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_48;
      7'b0110001 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_49;
      7'b0110010 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_50;
      7'b0110011 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_51;
      7'b0110100 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_52;
      7'b0110101 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_53;
      7'b0110110 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_54;
      7'b0110111 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_55;
      7'b0111000 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_56;
      7'b0111001 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_57;
      7'b0111010 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_58;
      7'b0111011 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_59;
      7'b0111100 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_60;
      7'b0111101 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_61;
      7'b0111110 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_62;
      7'b0111111 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_63;
      7'b1000000 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_64;
      7'b1000001 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_65;
      7'b1000010 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_66;
      7'b1000011 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_67;
      7'b1000100 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_68;
      7'b1000101 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_69;
      7'b1000110 : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_70;
      default : _zz__zz_when_PictureGenerator_l138_8_1 = fontVec_4_71;
    endcase
  end

  always @(*) begin
    case(_zz__zz_when_PictureGenerator_l138_8_10)
      7'b0000000 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_0;
      7'b0000001 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_1;
      7'b0000010 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_2;
      7'b0000011 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_3;
      7'b0000100 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_4;
      7'b0000101 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_5;
      7'b0000110 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_6;
      7'b0000111 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_7;
      7'b0001000 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_8;
      7'b0001001 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_9;
      7'b0001010 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_10;
      7'b0001011 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_11;
      7'b0001100 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_12;
      7'b0001101 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_13;
      7'b0001110 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_14;
      7'b0001111 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_15;
      7'b0010000 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_16;
      7'b0010001 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_17;
      7'b0010010 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_18;
      7'b0010011 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_19;
      7'b0010100 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_20;
      7'b0010101 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_21;
      7'b0010110 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_22;
      7'b0010111 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_23;
      7'b0011000 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_24;
      7'b0011001 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_25;
      7'b0011010 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_26;
      7'b0011011 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_27;
      7'b0011100 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_28;
      7'b0011101 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_29;
      7'b0011110 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_30;
      7'b0011111 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_31;
      7'b0100000 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_32;
      7'b0100001 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_33;
      7'b0100010 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_34;
      7'b0100011 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_35;
      7'b0100100 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_36;
      7'b0100101 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_37;
      7'b0100110 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_38;
      7'b0100111 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_39;
      7'b0101000 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_40;
      7'b0101001 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_41;
      7'b0101010 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_42;
      7'b0101011 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_43;
      7'b0101100 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_44;
      7'b0101101 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_45;
      7'b0101110 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_46;
      7'b0101111 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_47;
      7'b0110000 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_48;
      7'b0110001 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_49;
      7'b0110010 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_50;
      7'b0110011 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_51;
      7'b0110100 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_52;
      7'b0110101 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_53;
      7'b0110110 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_54;
      7'b0110111 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_55;
      7'b0111000 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_56;
      7'b0111001 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_57;
      7'b0111010 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_58;
      7'b0111011 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_59;
      7'b0111100 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_60;
      7'b0111101 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_61;
      7'b0111110 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_62;
      7'b0111111 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_63;
      7'b1000000 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_64;
      7'b1000001 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_65;
      7'b1000010 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_66;
      7'b1000011 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_67;
      7'b1000100 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_68;
      7'b1000101 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_69;
      7'b1000110 : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_70;
      default : _zz__zz_when_PictureGenerator_l138_8_9 = fontVec_4_71;
    endcase
  end

  always @(*) begin
    case(_zz__zz_when_PictureGenerator_l138_8_19)
      7'b0000000 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_0;
      7'b0000001 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_1;
      7'b0000010 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_2;
      7'b0000011 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_3;
      7'b0000100 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_4;
      7'b0000101 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_5;
      7'b0000110 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_6;
      7'b0000111 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_7;
      7'b0001000 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_8;
      7'b0001001 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_9;
      7'b0001010 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_10;
      7'b0001011 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_11;
      7'b0001100 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_12;
      7'b0001101 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_13;
      7'b0001110 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_14;
      7'b0001111 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_15;
      7'b0010000 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_16;
      7'b0010001 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_17;
      7'b0010010 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_18;
      7'b0010011 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_19;
      7'b0010100 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_20;
      7'b0010101 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_21;
      7'b0010110 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_22;
      7'b0010111 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_23;
      7'b0011000 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_24;
      7'b0011001 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_25;
      7'b0011010 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_26;
      7'b0011011 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_27;
      7'b0011100 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_28;
      7'b0011101 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_29;
      7'b0011110 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_30;
      7'b0011111 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_31;
      7'b0100000 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_32;
      7'b0100001 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_33;
      7'b0100010 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_34;
      7'b0100011 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_35;
      7'b0100100 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_36;
      7'b0100101 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_37;
      7'b0100110 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_38;
      7'b0100111 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_39;
      7'b0101000 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_40;
      7'b0101001 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_41;
      7'b0101010 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_42;
      7'b0101011 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_43;
      7'b0101100 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_44;
      7'b0101101 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_45;
      7'b0101110 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_46;
      7'b0101111 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_47;
      7'b0110000 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_48;
      7'b0110001 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_49;
      7'b0110010 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_50;
      7'b0110011 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_51;
      7'b0110100 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_52;
      7'b0110101 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_53;
      7'b0110110 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_54;
      7'b0110111 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_55;
      7'b0111000 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_56;
      7'b0111001 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_57;
      7'b0111010 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_58;
      7'b0111011 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_59;
      7'b0111100 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_60;
      7'b0111101 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_61;
      7'b0111110 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_62;
      7'b0111111 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_63;
      7'b1000000 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_64;
      7'b1000001 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_65;
      7'b1000010 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_66;
      7'b1000011 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_67;
      7'b1000100 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_68;
      7'b1000101 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_69;
      7'b1000110 : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_70;
      default : _zz__zz_when_PictureGenerator_l138_8_18 = fontVec_4_71;
    endcase
  end

  assign currXDiv = _zz_currXDiv;
  assign currYDiv = _zz_currYDiv;
  assign fontVec_0_0 = 8'h00;
  assign fontVec_0_1 = 8'h00;
  assign fontVec_0_2 = 8'h00;
  assign fontVec_0_3 = 8'h00;
  assign fontVec_0_4 = 8'h00;
  assign fontVec_0_5 = 8'h00;
  assign fontVec_0_6 = 8'h10;
  assign fontVec_0_7 = 8'h00;
  assign fontVec_0_8 = 8'h00;
  assign fontVec_0_9 = 8'h0c;
  assign fontVec_0_10 = 8'h7f;
  assign fontVec_0_11 = 8'hfc;
  assign fontVec_0_12 = 8'h04;
  assign fontVec_0_13 = 8'h40;
  assign fontVec_0_14 = 8'h08;
  assign fontVec_0_15 = 8'h04;
  assign fontVec_0_16 = 8'h40;
  assign fontVec_0_17 = 8'h08;
  assign fontVec_0_18 = 8'h00;
  assign fontVec_0_19 = 8'h40;
  assign fontVec_0_20 = 8'h08;
  assign fontVec_0_21 = 8'h41;
  assign fontVec_0_22 = 8'h5f;
  assign fontVec_0_23 = 8'he8;
  assign fontVec_0_24 = 8'h31;
  assign fontVec_0_25 = 8'h40;
  assign fontVec_0_26 = 8'h08;
  assign fontVec_0_27 = 8'h12;
  assign fontVec_0_28 = 8'h40;
  assign fontVec_0_29 = 8'h08;
  assign fontVec_0_30 = 8'h12;
  assign fontVec_0_31 = 8'h4f;
  assign fontVec_0_32 = 8'hc8;
  assign fontVec_0_33 = 8'h02;
  assign fontVec_0_34 = 8'h48;
  assign fontVec_0_35 = 8'h48;
  assign fontVec_0_36 = 8'h04;
  assign fontVec_0_37 = 8'h48;
  assign fontVec_0_38 = 8'h48;
  assign fontVec_0_39 = 8'h04;
  assign fontVec_0_40 = 8'h48;
  assign fontVec_0_41 = 8'h48;
  assign fontVec_0_42 = 8'h08;
  assign fontVec_0_43 = 8'h48;
  assign fontVec_0_44 = 8'h48;
  assign fontVec_0_45 = 8'h08;
  assign fontVec_0_46 = 8'h4f;
  assign fontVec_0_47 = 8'hc8;
  assign fontVec_0_48 = 8'h38;
  assign fontVec_0_49 = 8'h48;
  assign fontVec_0_50 = 8'h48;
  assign fontVec_0_51 = 8'h18;
  assign fontVec_0_52 = 8'h48;
  assign fontVec_0_53 = 8'h08;
  assign fontVec_0_54 = 8'h18;
  assign fontVec_0_55 = 8'h40;
  assign fontVec_0_56 = 8'h08;
  assign fontVec_0_57 = 8'h18;
  assign fontVec_0_58 = 8'h40;
  assign fontVec_0_59 = 8'h08;
  assign fontVec_0_60 = 8'h18;
  assign fontVec_0_61 = 8'h40;
  assign fontVec_0_62 = 8'h08;
  assign fontVec_0_63 = 8'h00;
  assign fontVec_0_64 = 8'h40;
  assign fontVec_0_65 = 8'h38;
  assign fontVec_0_66 = 8'h00;
  assign fontVec_0_67 = 8'h40;
  assign fontVec_0_68 = 8'h18;
  assign fontVec_0_69 = 8'h00;
  assign fontVec_0_70 = 8'h00;
  assign fontVec_0_71 = 8'h00;
  assign fontVec_1_0 = 8'h00;
  assign fontVec_1_1 = 8'h00;
  assign fontVec_1_2 = 8'h00;
  assign fontVec_1_3 = 8'h00;
  assign fontVec_1_4 = 8'h10;
  assign fontVec_1_5 = 8'h00;
  assign fontVec_1_6 = 8'h00;
  assign fontVec_1_7 = 8'h08;
  assign fontVec_1_8 = 8'h00;
  assign fontVec_1_9 = 8'h00;
  assign fontVec_1_10 = 8'h08;
  assign fontVec_1_11 = 8'h00;
  assign fontVec_1_12 = 8'h0f;
  assign fontVec_1_13 = 8'hff;
  assign fontVec_1_14 = 8'hfc;
  assign fontVec_1_15 = 8'h11;
  assign fontVec_1_16 = 8'h00;
  assign fontVec_1_17 = 8'h08;
  assign fontVec_1_18 = 8'h33;
  assign fontVec_1_19 = 8'h04;
  assign fontVec_1_20 = 8'h10;
  assign fontVec_1_21 = 8'h03;
  assign fontVec_1_22 = 8'hff;
  assign fontVec_1_23 = 8'hf8;
  assign fontVec_1_24 = 8'h04;
  assign fontVec_1_25 = 8'h32;
  assign fontVec_1_26 = 8'h10;
  assign fontVec_1_27 = 8'h0f;
  assign fontVec_1_28 = 8'h22;
  assign fontVec_1_29 = 8'h20;
  assign fontVec_1_30 = 8'h09;
  assign fontVec_1_31 = 8'h41;
  assign fontVec_1_32 = 8'h40;
  assign fontVec_1_33 = 8'h19;
  assign fontVec_1_34 = 8'hc3;
  assign fontVec_1_35 = 8'h80;
  assign fontVec_1_36 = 8'h24;
  assign fontVec_1_37 = 8'hff;
  assign fontVec_1_38 = 8'hc0;
  assign fontVec_1_39 = 8'h07;
  assign fontVec_1_40 = 8'h00;
  assign fontVec_1_41 = 8'h70;
  assign fontVec_1_42 = 8'h04;
  assign fontVec_1_43 = 8'h00;
  assign fontVec_1_44 = 8'h5e;
  assign fontVec_1_45 = 8'h1f;
  assign fontVec_1_46 = 8'hff;
  assign fontVec_1_47 = 8'he8;
  assign fontVec_1_48 = 8'h20;
  assign fontVec_1_49 = 8'h18;
  assign fontVec_1_50 = 8'h10;
  assign fontVec_1_51 = 8'h01;
  assign fontVec_1_52 = 8'h99;
  assign fontVec_1_53 = 8'h00;
  assign fontVec_1_54 = 8'h03;
  assign fontVec_1_55 = 8'h18;
  assign fontVec_1_56 = 8'h80;
  assign fontVec_1_57 = 8'h06;
  assign fontVec_1_58 = 8'h18;
  assign fontVec_1_59 = 8'h60;
  assign fontVec_1_60 = 8'h08;
  assign fontVec_1_61 = 8'h18;
  assign fontVec_1_62 = 8'h30;
  assign fontVec_1_63 = 8'h10;
  assign fontVec_1_64 = 8'h78;
  assign fontVec_1_65 = 8'h10;
  assign fontVec_1_66 = 8'h00;
  assign fontVec_1_67 = 8'h10;
  assign fontVec_1_68 = 8'h00;
  assign fontVec_1_69 = 8'h00;
  assign fontVec_1_70 = 8'h00;
  assign fontVec_1_71 = 8'h00;
  assign fontVec_2_0 = 8'h00;
  assign fontVec_2_1 = 8'h00;
  assign fontVec_2_2 = 8'h00;
  assign fontVec_2_3 = 8'h00;
  assign fontVec_2_4 = 8'h00;
  assign fontVec_2_5 = 8'h30;
  assign fontVec_2_6 = 8'h00;
  assign fontVec_2_7 = 8'h03;
  assign fontVec_2_8 = 8'hf8;
  assign fontVec_2_9 = 8'h3f;
  assign fontVec_2_10 = 8'h7c;
  assign fontVec_2_11 = 8'h00;
  assign fontVec_2_12 = 8'h22;
  assign fontVec_2_13 = 8'h20;
  assign fontVec_2_14 = 8'h10;
  assign fontVec_2_15 = 8'h22;
  assign fontVec_2_16 = 8'h32;
  assign fontVec_2_17 = 8'h30;
  assign fontVec_2_18 = 8'h22;
  assign fontVec_2_19 = 8'h13;
  assign fontVec_2_20 = 8'h20;
  assign fontVec_2_21 = 8'h22;
  assign fontVec_2_22 = 8'h12;
  assign fontVec_2_23 = 8'h40;
  assign fontVec_2_24 = 8'h3e;
  assign fontVec_2_25 = 8'h7f;
  assign fontVec_2_26 = 8'hfc;
  assign fontVec_2_27 = 8'h22;
  assign fontVec_2_28 = 8'h40;
  assign fontVec_2_29 = 8'h0c;
  assign fontVec_2_30 = 8'h22;
  assign fontVec_2_31 = 8'hf0;
  assign fontVec_2_32 = 8'h38;
  assign fontVec_2_33 = 8'h22;
  assign fontVec_2_34 = 8'h20;
  assign fontVec_2_35 = 8'h28;
  assign fontVec_2_36 = 8'h22;
  assign fontVec_2_37 = 8'h3f;
  assign fontVec_2_38 = 8'hfc;
  assign fontVec_2_39 = 8'h3e;
  assign fontVec_2_40 = 8'h4d;
  assign fontVec_2_41 = 8'h20;
  assign fontVec_2_42 = 8'h22;
  assign fontVec_2_43 = 8'h89;
  assign fontVec_2_44 = 8'h20;
  assign fontVec_2_45 = 8'h23;
  assign fontVec_2_46 = 8'heb;
  assign fontVec_2_47 = 8'h20;
  assign fontVec_2_48 = 8'h22;
  assign fontVec_2_49 = 8'h33;
  assign fontVec_2_50 = 8'hfc;
  assign fontVec_2_51 = 8'h22;
  assign fontVec_2_52 = 8'h10;
  assign fontVec_2_53 = 8'h20;
  assign fontVec_2_54 = 8'h3e;
  assign fontVec_2_55 = 8'h20;
  assign fontVec_2_56 = 8'h20;
  assign fontVec_2_57 = 8'h22;
  assign fontVec_2_58 = 8'h40;
  assign fontVec_2_59 = 8'h20;
  assign fontVec_2_60 = 8'h20;
  assign fontVec_2_61 = 8'h80;
  assign fontVec_2_62 = 8'h20;
  assign fontVec_2_63 = 8'h23;
  assign fontVec_2_64 = 8'h00;
  assign fontVec_2_65 = 8'h20;
  assign fontVec_2_66 = 8'h04;
  assign fontVec_2_67 = 8'h00;
  assign fontVec_2_68 = 8'h20;
  assign fontVec_2_69 = 8'h00;
  assign fontVec_2_70 = 8'h00;
  assign fontVec_2_71 = 8'h00;
  assign fontVec_3_0 = 8'h00;
  assign fontVec_3_1 = 8'h00;
  assign fontVec_3_2 = 8'h00;
  assign fontVec_3_3 = 8'h00;
  assign fontVec_3_4 = 8'h30;
  assign fontVec_3_5 = 8'h00;
  assign fontVec_3_6 = 8'h00;
  assign fontVec_3_7 = 8'h20;
  assign fontVec_3_8 = 8'h00;
  assign fontVec_3_9 = 8'h03;
  assign fontVec_3_10 = 8'hff;
  assign fontVec_3_11 = 8'he0;
  assign fontVec_3_12 = 8'h02;
  assign fontVec_3_13 = 8'h00;
  assign fontVec_3_14 = 8'h40;
  assign fontVec_3_15 = 8'h02;
  assign fontVec_3_16 = 8'h00;
  assign fontVec_3_17 = 8'h40;
  assign fontVec_3_18 = 8'h03;
  assign fontVec_3_19 = 8'hff;
  assign fontVec_3_20 = 8'hc0;
  assign fontVec_3_21 = 8'h02;
  assign fontVec_3_22 = 8'h00;
  assign fontVec_3_23 = 8'h40;
  assign fontVec_3_24 = 8'h02;
  assign fontVec_3_25 = 8'h00;
  assign fontVec_3_26 = 8'h40;
  assign fontVec_3_27 = 8'h03;
  assign fontVec_3_28 = 8'hff;
  assign fontVec_3_29 = 8'hc0;
  assign fontVec_3_30 = 8'h02;
  assign fontVec_3_31 = 8'h00;
  assign fontVec_3_32 = 8'h40;
  assign fontVec_3_33 = 8'h02;
  assign fontVec_3_34 = 8'h00;
  assign fontVec_3_35 = 8'h40;
  assign fontVec_3_36 = 8'h03;
  assign fontVec_3_37 = 8'hff;
  assign fontVec_3_38 = 8'he0;
  assign fontVec_3_39 = 8'h02;
  assign fontVec_3_40 = 8'h20;
  assign fontVec_3_41 = 8'h40;
  assign fontVec_3_42 = 8'h00;
  assign fontVec_3_43 = 8'h10;
  assign fontVec_3_44 = 8'h00;
  assign fontVec_3_45 = 8'h01;
  assign fontVec_3_46 = 8'h18;
  assign fontVec_3_47 = 8'h00;
  assign fontVec_3_48 = 8'h09;
  assign fontVec_3_49 = 8'h8c;
  assign fontVec_3_50 = 8'h10;
  assign fontVec_3_51 = 8'h09;
  assign fontVec_3_52 = 8'h8c;
  assign fontVec_3_53 = 8'h08;
  assign fontVec_3_54 = 8'h09;
  assign fontVec_3_55 = 8'h80;
  assign fontVec_3_56 = 8'h4c;
  assign fontVec_3_57 = 8'h19;
  assign fontVec_3_58 = 8'h80;
  assign fontVec_3_59 = 8'h44;
  assign fontVec_3_60 = 8'h38;
  assign fontVec_3_61 = 8'h80;
  assign fontVec_3_62 = 8'hc4;
  assign fontVec_3_63 = 8'h00;
  assign fontVec_3_64 = 8'hff;
  assign fontVec_3_65 = 8'hc0;
  assign fontVec_3_66 = 8'h00;
  assign fontVec_3_67 = 8'h00;
  assign fontVec_3_68 = 8'h00;
  assign fontVec_3_69 = 8'h00;
  assign fontVec_3_70 = 8'h00;
  assign fontVec_3_71 = 8'h00;
  assign fontVec_4_0 = 8'h00;
  assign fontVec_4_1 = 8'h00;
  assign fontVec_4_2 = 8'h00;
  assign fontVec_4_3 = 8'h00;
  assign fontVec_4_4 = 8'h00;
  assign fontVec_4_5 = 8'h00;
  assign fontVec_4_6 = 8'h00;
  assign fontVec_4_7 = 8'h02;
  assign fontVec_4_8 = 8'h00;
  assign fontVec_4_9 = 8'h1f;
  assign fontVec_4_10 = 8'hc3;
  assign fontVec_4_11 = 8'h00;
  assign fontVec_4_12 = 8'h10;
  assign fontVec_4_13 = 8'hc3;
  assign fontVec_4_14 = 8'h00;
  assign fontVec_4_15 = 8'h10;
  assign fontVec_4_16 = 8'h83;
  assign fontVec_4_17 = 8'h00;
  assign fontVec_4_18 = 8'h10;
  assign fontVec_4_19 = 8'h83;
  assign fontVec_4_20 = 8'h00;
  assign fontVec_4_21 = 8'h11;
  assign fontVec_4_22 = 8'h03;
  assign fontVec_4_23 = 8'h00;
  assign fontVec_4_24 = 8'h11;
  assign fontVec_4_25 = 8'h03;
  assign fontVec_4_26 = 8'h00;
  assign fontVec_4_27 = 8'h12;
  assign fontVec_4_28 = 8'h03;
  assign fontVec_4_29 = 8'h00;
  assign fontVec_4_30 = 8'h12;
  assign fontVec_4_31 = 8'h02;
  assign fontVec_4_32 = 8'h80;
  assign fontVec_4_33 = 8'h11;
  assign fontVec_4_34 = 8'h02;
  assign fontVec_4_35 = 8'h80;
  assign fontVec_4_36 = 8'h10;
  assign fontVec_4_37 = 8'h86;
  assign fontVec_4_38 = 8'h80;
  assign fontVec_4_39 = 8'h10;
  assign fontVec_4_40 = 8'hc4;
  assign fontVec_4_41 = 8'h80;
  assign fontVec_4_42 = 8'h10;
  assign fontVec_4_43 = 8'h44;
  assign fontVec_4_44 = 8'h80;
  assign fontVec_4_45 = 8'h10;
  assign fontVec_4_46 = 8'h44;
  assign fontVec_4_47 = 8'h40;
  assign fontVec_4_48 = 8'h10;
  assign fontVec_4_49 = 8'h48;
  assign fontVec_4_50 = 8'h40;
  assign fontVec_4_51 = 8'h17;
  assign fontVec_4_52 = 8'hc8;
  assign fontVec_4_53 = 8'h60;
  assign fontVec_4_54 = 8'h11;
  assign fontVec_4_55 = 8'h90;
  assign fontVec_4_56 = 8'h20;
  assign fontVec_4_57 = 8'h10;
  assign fontVec_4_58 = 8'h30;
  assign fontVec_4_59 = 8'h30;
  assign fontVec_4_60 = 8'h10;
  assign fontVec_4_61 = 8'h60;
  assign fontVec_4_62 = 8'h18;
  assign fontVec_4_63 = 8'h10;
  assign fontVec_4_64 = 8'h80;
  assign fontVec_4_65 = 8'h0e;
  assign fontVec_4_66 = 8'h11;
  assign fontVec_4_67 = 8'h00;
  assign fontVec_4_68 = 8'h00;
  assign fontVec_4_69 = 8'h00;
  assign fontVec_4_70 = 8'h00;
  assign fontVec_4_71 = 8'h00;
  always @(*) begin
    color_rgb = 16'h0000;
    if(when_PictureGenerator_l97) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_1) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_2) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_3) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_4) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_5) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_6) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_7) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_8) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_9) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_10) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_11) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_12) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_13) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_14) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_15) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_16) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_17) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_18) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_19) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_20) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_21) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_22) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_23) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_24) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_25) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_26) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_27) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_28) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_29) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_30) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_31) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_32) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_33) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_34) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_35) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_36) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_37) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_38) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_39) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_40) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_41) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_42) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_43) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_44) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_45) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_46) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_47) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_48) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_49) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_50) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_51) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_52) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_53) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_54) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_55) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_56) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_57) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_58) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_59) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_60) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_61) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_62) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_63) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_64) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_65) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_66) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_67) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_68) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_69) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_70) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_71) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_72) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_73) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_74) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_75) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_76) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_77) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_78) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_79) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_80) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_81) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_82) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_83) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_84) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_85) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_86) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_87) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_88) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_89) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_90) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_91) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_92) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_93) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_94) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_95) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_96) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_97) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_98) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_99) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_100) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_101) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_102) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_103) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_104) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_105) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_106) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_107) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_108) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_109) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_110) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_111) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_112) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_113) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_114) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_115) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_116) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_117) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_118) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_119) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_120) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_121) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_122) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_123) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_124) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_125) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_126) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_127) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_128) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_129) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_130) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_131) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_132) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_133) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_134) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_135) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_136) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_137) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_138) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_139) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_140) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_141) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_142) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_143) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_144) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_145) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_146) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_147) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_148) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_149) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_150) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_151) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_152) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_153) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_154) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_155) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_156) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_157) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_158) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_159) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_160) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_161) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_162) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_163) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_164) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_165) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_166) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_167) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_168) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_169) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_170) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_171) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_172) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_173) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_174) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_175) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_176) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_177) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_178) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_179) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_180) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_181) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_182) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_183) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_184) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_185) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_186) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_187) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_188) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_189) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_190) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_191) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_192) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_193) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_194) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_195) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_196) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_197) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_198) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_199) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_200) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_201) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_202) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_203) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_204) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_205) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_206) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_207) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_208) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_209) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_210) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_211) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_212) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_213) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_214) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_215) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_216) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_217) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_218) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_219) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_220) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_221) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_222) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_223) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_224) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_225) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_226) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_227) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_228) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_229) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_230) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_231) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_232) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_233) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_234) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_235) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_236) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_237) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_238) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_239) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_240) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_241) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_242) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_243) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_244) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_245) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_246) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_247) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_248) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_249) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_250) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_251) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_252) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_253) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_254) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_255) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_256) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_257) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_258) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_259) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_260) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_261) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_262) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_263) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_264) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_265) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_266) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_267) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_268) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_269) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_270) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_271) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_272) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_273) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_274) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_275) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_276) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_277) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_278) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_279) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_280) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_281) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_282) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_283) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_284) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_285) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_286) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_287) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_288) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_289) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_290) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_291) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_292) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_293) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_294) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_295) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_296) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_297) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_298) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_299) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_300) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_301) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_302) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_303) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_304) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_305) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_306) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_307) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_308) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_309) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_310) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_311) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_312) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_313) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_314) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_315) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_316) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_317) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_318) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_319) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_320) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_321) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_322) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_323) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_324) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_325) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_326) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_327) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_328) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_329) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_330) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_331) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_332) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_333) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_334) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_335) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_336) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_337) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_338) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_339) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_340) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_341) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_342) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_343) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_344) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_345) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_346) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_347) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_348) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_349) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_350) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_351) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_352) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_353) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_354) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_355) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_356) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_357) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_358) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_359) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_360) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_361) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_362) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_363) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_364) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_365) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_366) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_367) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_368) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_369) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_370) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_371) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_372) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_373) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_374) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_375) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_376) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_377) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_378) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_379) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_380) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_381) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_382) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_383) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_384) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_385) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_386) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_387) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_388) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_389) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_390) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_391) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_392) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_393) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_394) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_395) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_396) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_397) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_398) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_399) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_400) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_401) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_402) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_403) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_404) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_405) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_406) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_407) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_408) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_409) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_410) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_411) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_412) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_413) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_414) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_415) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_416) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_417) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_418) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_419) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_420) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_421) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_422) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_423) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_424) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_425) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_426) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_427) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_428) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_429) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_430) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_431) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_432) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_433) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_434) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_435) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_436) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_437) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_438) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_439) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_440) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_441) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_442) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_443) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_444) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_445) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_446) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_447) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_448) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_449) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_450) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_451) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_452) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_453) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_454) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_455) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_456) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_457) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_458) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_459) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_460) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_461) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_462) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_463) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_464) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_465) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_466) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_467) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_468) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_469) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_470) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_471) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_472) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_473) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_474) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_475) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_476) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_477) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_478) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_479) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_480) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_481) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_482) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_483) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_484) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_485) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_486) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_487) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_488) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_489) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_490) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_491) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_492) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_493) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_494) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_495) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_496) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_497) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_498) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_499) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_500) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_501) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_502) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_503) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_504) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_505) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_506) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_507) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_508) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_509) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_510) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_511) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_512) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_513) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_514) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_515) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_516) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_517) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_518) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_519) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_520) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_521) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_522) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_523) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_524) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_525) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_526) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_527) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_528) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_529) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_530) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_531) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_532) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_533) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_534) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_535) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_536) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_537) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_538) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_539) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_540) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_541) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_542) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_543) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_544) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_545) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_546) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_547) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_548) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_549) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_550) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_551) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_552) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_553) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_554) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_555) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_556) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_557) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_558) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_559) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_560) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_561) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_562) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_563) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_564) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_565) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_566) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_567) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_568) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_569) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_570) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_571) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_572) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_573) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_574) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_575) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_576) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_577) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_578) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_579) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_580) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_581) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_582) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_583) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_584) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_585) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_586) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_587) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_588) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_589) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_590) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_591) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_592) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_593) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_594) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_595) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_596) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_597) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_598) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_599) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_600) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_601) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_602) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_603) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_604) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_605) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_606) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_607) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_608) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_609) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_610) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_611) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_612) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_613) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_614) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_615) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_616) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_617) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_618) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_619) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_620) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_621) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_622) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_623) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_624) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_625) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_626) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_627) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_628) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l102_629) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_1) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_2) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_3) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_4) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_5) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_6) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_7) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_8) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_9) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_10) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_11) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_12) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_13) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_14) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_15) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_16) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_17) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_18) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_19) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_20) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_21) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_22) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_23) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_24) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_25) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_26) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_27) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_28) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_29) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_30) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_31) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_32) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_33) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_34) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_35) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_36) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_37) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_38) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_39) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_40) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_41) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_42) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_43) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_44) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_45) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_46) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_47) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_48) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_49) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_50) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_51) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_52) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_53) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_54) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_55) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_56) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_57) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_58) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_59) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_60) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_61) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_62) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_63) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_64) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_65) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_66) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_67) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_68) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_69) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_70) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_71) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_72) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_73) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_74) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_75) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_76) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_77) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_78) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_79) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_80) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_81) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_82) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_83) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_84) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_85) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_86) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_87) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_88) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_89) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_90) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_91) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_92) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_93) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_94) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_95) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_96) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_97) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_98) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_99) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_100) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_101) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_102) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_103) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_104) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_105) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_106) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_107) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_108) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_109) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_110) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_111) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_112) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_113) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_114) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_115) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_116) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_117) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_118) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_119) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_120) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_121) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_122) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_123) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_124) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_125) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_126) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_127) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_128) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_129) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_130) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_131) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_132) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_133) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_134) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_135) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_136) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_137) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_138) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_139) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_140) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_141) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_142) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_143) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_144) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_145) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_146) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_147) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_148) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_149) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_150) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_151) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_152) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_153) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_154) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_155) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_156) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_157) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_158) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_159) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_160) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_161) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_162) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_163) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_164) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_165) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_166) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_167) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_168) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_169) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_170) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_171) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_172) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_173) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_174) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_175) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_176) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_177) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_178) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_179) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_180) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_181) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_182) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_183) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_184) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_185) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_186) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_187) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_188) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_189) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_190) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_191) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_192) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_193) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_194) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_195) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_196) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_197) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_198) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_199) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_200) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_201) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_202) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_203) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_204) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_205) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_206) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_207) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_208) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_209) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_210) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_211) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_212) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_213) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_214) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_215) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_216) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_217) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_218) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_219) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_220) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_221) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_222) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_223) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_224) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_225) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_226) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_227) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_228) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_229) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_230) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_231) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_232) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_233) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_234) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_235) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_236) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_237) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_238) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_239) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_240) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_241) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_242) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_243) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_244) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_245) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_246) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_247) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_248) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_249) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_250) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_251) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_252) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_253) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_254) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_255) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_256) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_257) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_258) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_259) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_260) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_261) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_262) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_263) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_264) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_265) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_266) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_267) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_268) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_269) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_270) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_271) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_272) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_273) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_274) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_275) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_276) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_277) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_278) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_279) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_280) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_281) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_282) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_283) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_284) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_285) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_286) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_287) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_288) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_289) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_290) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_291) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_292) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_293) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_294) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_295) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_296) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_297) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_298) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_299) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_300) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_301) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_302) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_303) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_304) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_305) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_306) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_307) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_308) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_309) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_310) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_311) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_312) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_313) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_314) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_315) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_316) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_317) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_318) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_319) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_320) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_321) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_322) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_323) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_324) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_325) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_326) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_327) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_328) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_329) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_330) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_331) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_332) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_333) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_334) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_335) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_336) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_337) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_338) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_339) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_340) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_341) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_342) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_343) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_344) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_345) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_346) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_347) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_348) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_349) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_350) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_351) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_352) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_353) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_354) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_355) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_356) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_357) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_358) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_359) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_360) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_361) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_362) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_363) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_364) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_365) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_366) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_367) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_368) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_369) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_370) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_371) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_372) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_373) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_374) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_375) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_376) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_377) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_378) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_379) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_380) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_381) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_382) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_383) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_384) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_385) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_386) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_387) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_388) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_389) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_390) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_391) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_392) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_393) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_394) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_395) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_396) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_397) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_398) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_399) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_400) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_401) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_402) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_403) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_404) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_405) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_406) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_407) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_408) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_409) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_410) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_411) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_412) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_413) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_414) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_415) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_416) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_417) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_418) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_419) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_420) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_421) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_422) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_423) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_424) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_425) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_426) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_427) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_428) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_429) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_430) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_431) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_432) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_433) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_434) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_435) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_436) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_437) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_438) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_439) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_440) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_441) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_442) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_443) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_444) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_445) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_446) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_447) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_448) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_449) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_450) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_451) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_452) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_453) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_454) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_455) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_456) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_457) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_458) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_459) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_460) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_461) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_462) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_463) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_464) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_465) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_466) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_467) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_468) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_469) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_470) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_471) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_472) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_473) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_474) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_475) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_476) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_477) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_478) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_479) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_480) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_481) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_482) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_483) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_484) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_485) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_486) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_487) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_488) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_489) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_490) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_491) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_492) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_493) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_494) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_495) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_496) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_497) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_498) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_499) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_500) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_501) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_502) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_503) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_504) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_505) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_506) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_507) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_508) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_509) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_510) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_511) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_512) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_513) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_514) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_515) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_516) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l110_517) begin
      color_rgb = 16'h6b4d;
    end
    if(when_PictureGenerator_l115) begin
      color_rgb = 16'hffff;
    end else begin
      if(when_PictureGenerator_l117) begin
        color_rgb = 16'hffff;
      end else begin
        if(when_PictureGenerator_l119) begin
          color_rgb = colorInRam;
        end else begin
          if(when_PictureGenerator_l121) begin
            color_rgb = 16'h6b4d;
          end
        end
      end
    end
    if(when_PictureGenerator_l138) begin
      color_rgb = 16'hffff;
    end
    if(when_PictureGenerator_l138_1) begin
      color_rgb = 16'hffff;
    end
    if(when_PictureGenerator_l138_2) begin
      color_rgb = 16'hffff;
    end
    if(when_PictureGenerator_l138_3) begin
      color_rgb = 16'hffff;
    end
    if(when_PictureGenerator_l138_4) begin
      color_rgb = 16'hffff;
    end
  end

  assign when_PictureGenerator_l97 = (((10'h027 < currYDiv) && (currYDiv < 10'h129)) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102 = ((currYDiv == 10'h02c) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_1 = ((currYDiv == 10'h030) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_2 = ((currYDiv == 10'h034) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_3 = ((currYDiv == 10'h038) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_4 = ((currYDiv == 10'h03c) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_5 = ((currYDiv == 10'h040) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_6 = ((currYDiv == 10'h044) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_7 = ((currYDiv == 10'h048) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_8 = ((currYDiv == 10'h04c) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_9 = ((currYDiv == 10'h050) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_10 = ((currYDiv == 10'h054) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_11 = ((currYDiv == 10'h058) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_12 = ((currYDiv == 10'h05c) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_13 = ((currYDiv == 10'h060) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_14 = ((currYDiv == 10'h064) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_15 = ((currYDiv == 10'h068) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_16 = ((currYDiv == 10'h06c) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_17 = ((currYDiv == 10'h070) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_18 = ((currYDiv == 10'h074) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_19 = ((currYDiv == 10'h078) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_20 = ((currYDiv == 10'h07c) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_21 = ((currYDiv == 10'h080) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_22 = ((currYDiv == 10'h084) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_23 = ((currYDiv == 10'h088) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_24 = ((currYDiv == 10'h08c) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_25 = ((currYDiv == 10'h090) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_26 = ((currYDiv == 10'h094) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_27 = ((currYDiv == 10'h098) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_28 = ((currYDiv == 10'h09c) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_29 = ((currYDiv == 10'h0a0) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_30 = ((currYDiv == 10'h0a4) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_31 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_32 = ((currYDiv == 10'h0ac) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_33 = ((currYDiv == 10'h0b0) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_34 = ((currYDiv == 10'h0b4) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_35 = ((currYDiv == 10'h0b8) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_36 = ((currYDiv == 10'h0bc) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_37 = ((currYDiv == 10'h0c0) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_38 = ((currYDiv == 10'h0c4) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_39 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_40 = ((currYDiv == 10'h0cc) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_41 = ((currYDiv == 10'h0d0) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_42 = ((currYDiv == 10'h0d4) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_43 = ((currYDiv == 10'h0d8) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_44 = ((currYDiv == 10'h0dc) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_45 = ((currYDiv == 10'h0e0) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_46 = ((currYDiv == 10'h0e4) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_47 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_48 = ((currYDiv == 10'h0ec) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_49 = ((currYDiv == 10'h0f0) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_50 = ((currYDiv == 10'h0f4) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_51 = ((currYDiv == 10'h0f8) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_52 = ((currYDiv == 10'h0fc) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_53 = ((currYDiv == 10'h100) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_54 = ((currYDiv == 10'h104) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_55 = ((currYDiv == 10'h108) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_56 = ((currYDiv == 10'h10c) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_57 = ((currYDiv == 10'h110) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_58 = ((currYDiv == 10'h114) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_59 = ((currYDiv == 10'h118) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_60 = ((currYDiv == 10'h11c) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_61 = ((currYDiv == 10'h120) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_62 = ((currYDiv == 10'h124) && (currXDiv == 10'h085));
  assign when_PictureGenerator_l102_63 = ((currYDiv == 10'h02c) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_64 = ((currYDiv == 10'h030) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_65 = ((currYDiv == 10'h034) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_66 = ((currYDiv == 10'h038) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_67 = ((currYDiv == 10'h03c) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_68 = ((currYDiv == 10'h040) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_69 = ((currYDiv == 10'h044) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_70 = ((currYDiv == 10'h048) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_71 = ((currYDiv == 10'h04c) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_72 = ((currYDiv == 10'h050) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_73 = ((currYDiv == 10'h054) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_74 = ((currYDiv == 10'h058) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_75 = ((currYDiv == 10'h05c) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_76 = ((currYDiv == 10'h060) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_77 = ((currYDiv == 10'h064) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_78 = ((currYDiv == 10'h068) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_79 = ((currYDiv == 10'h06c) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_80 = ((currYDiv == 10'h070) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_81 = ((currYDiv == 10'h074) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_82 = ((currYDiv == 10'h078) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_83 = ((currYDiv == 10'h07c) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_84 = ((currYDiv == 10'h080) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_85 = ((currYDiv == 10'h084) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_86 = ((currYDiv == 10'h088) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_87 = ((currYDiv == 10'h08c) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_88 = ((currYDiv == 10'h090) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_89 = ((currYDiv == 10'h094) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_90 = ((currYDiv == 10'h098) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_91 = ((currYDiv == 10'h09c) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_92 = ((currYDiv == 10'h0a0) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_93 = ((currYDiv == 10'h0a4) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_94 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_95 = ((currYDiv == 10'h0ac) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_96 = ((currYDiv == 10'h0b0) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_97 = ((currYDiv == 10'h0b4) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_98 = ((currYDiv == 10'h0b8) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_99 = ((currYDiv == 10'h0bc) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_100 = ((currYDiv == 10'h0c0) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_101 = ((currYDiv == 10'h0c4) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_102 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_103 = ((currYDiv == 10'h0cc) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_104 = ((currYDiv == 10'h0d0) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_105 = ((currYDiv == 10'h0d4) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_106 = ((currYDiv == 10'h0d8) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_107 = ((currYDiv == 10'h0dc) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_108 = ((currYDiv == 10'h0e0) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_109 = ((currYDiv == 10'h0e4) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_110 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_111 = ((currYDiv == 10'h0ec) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_112 = ((currYDiv == 10'h0f0) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_113 = ((currYDiv == 10'h0f4) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_114 = ((currYDiv == 10'h0f8) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_115 = ((currYDiv == 10'h0fc) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_116 = ((currYDiv == 10'h100) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_117 = ((currYDiv == 10'h104) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_118 = ((currYDiv == 10'h108) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_119 = ((currYDiv == 10'h10c) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_120 = ((currYDiv == 10'h110) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_121 = ((currYDiv == 10'h114) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_122 = ((currYDiv == 10'h118) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_123 = ((currYDiv == 10'h11c) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_124 = ((currYDiv == 10'h120) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_125 = ((currYDiv == 10'h124) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l102_126 = ((currYDiv == 10'h02c) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_127 = ((currYDiv == 10'h030) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_128 = ((currYDiv == 10'h034) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_129 = ((currYDiv == 10'h038) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_130 = ((currYDiv == 10'h03c) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_131 = ((currYDiv == 10'h040) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_132 = ((currYDiv == 10'h044) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_133 = ((currYDiv == 10'h048) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_134 = ((currYDiv == 10'h04c) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_135 = ((currYDiv == 10'h050) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_136 = ((currYDiv == 10'h054) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_137 = ((currYDiv == 10'h058) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_138 = ((currYDiv == 10'h05c) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_139 = ((currYDiv == 10'h060) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_140 = ((currYDiv == 10'h064) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_141 = ((currYDiv == 10'h068) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_142 = ((currYDiv == 10'h06c) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_143 = ((currYDiv == 10'h070) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_144 = ((currYDiv == 10'h074) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_145 = ((currYDiv == 10'h078) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_146 = ((currYDiv == 10'h07c) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_147 = ((currYDiv == 10'h080) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_148 = ((currYDiv == 10'h084) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_149 = ((currYDiv == 10'h088) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_150 = ((currYDiv == 10'h08c) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_151 = ((currYDiv == 10'h090) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_152 = ((currYDiv == 10'h094) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_153 = ((currYDiv == 10'h098) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_154 = ((currYDiv == 10'h09c) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_155 = ((currYDiv == 10'h0a0) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_156 = ((currYDiv == 10'h0a4) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_157 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_158 = ((currYDiv == 10'h0ac) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_159 = ((currYDiv == 10'h0b0) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_160 = ((currYDiv == 10'h0b4) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_161 = ((currYDiv == 10'h0b8) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_162 = ((currYDiv == 10'h0bc) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_163 = ((currYDiv == 10'h0c0) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_164 = ((currYDiv == 10'h0c4) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_165 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_166 = ((currYDiv == 10'h0cc) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_167 = ((currYDiv == 10'h0d0) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_168 = ((currYDiv == 10'h0d4) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_169 = ((currYDiv == 10'h0d8) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_170 = ((currYDiv == 10'h0dc) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_171 = ((currYDiv == 10'h0e0) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_172 = ((currYDiv == 10'h0e4) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_173 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_174 = ((currYDiv == 10'h0ec) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_175 = ((currYDiv == 10'h0f0) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_176 = ((currYDiv == 10'h0f4) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_177 = ((currYDiv == 10'h0f8) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_178 = ((currYDiv == 10'h0fc) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_179 = ((currYDiv == 10'h100) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_180 = ((currYDiv == 10'h104) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_181 = ((currYDiv == 10'h108) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_182 = ((currYDiv == 10'h10c) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_183 = ((currYDiv == 10'h110) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_184 = ((currYDiv == 10'h114) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_185 = ((currYDiv == 10'h118) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_186 = ((currYDiv == 10'h11c) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_187 = ((currYDiv == 10'h120) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_188 = ((currYDiv == 10'h124) && (currXDiv == 10'h0c1));
  assign when_PictureGenerator_l102_189 = ((currYDiv == 10'h02c) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_190 = ((currYDiv == 10'h030) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_191 = ((currYDiv == 10'h034) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_192 = ((currYDiv == 10'h038) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_193 = ((currYDiv == 10'h03c) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_194 = ((currYDiv == 10'h040) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_195 = ((currYDiv == 10'h044) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_196 = ((currYDiv == 10'h048) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_197 = ((currYDiv == 10'h04c) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_198 = ((currYDiv == 10'h050) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_199 = ((currYDiv == 10'h054) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_200 = ((currYDiv == 10'h058) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_201 = ((currYDiv == 10'h05c) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_202 = ((currYDiv == 10'h060) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_203 = ((currYDiv == 10'h064) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_204 = ((currYDiv == 10'h068) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_205 = ((currYDiv == 10'h06c) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_206 = ((currYDiv == 10'h070) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_207 = ((currYDiv == 10'h074) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_208 = ((currYDiv == 10'h078) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_209 = ((currYDiv == 10'h07c) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_210 = ((currYDiv == 10'h080) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_211 = ((currYDiv == 10'h084) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_212 = ((currYDiv == 10'h088) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_213 = ((currYDiv == 10'h08c) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_214 = ((currYDiv == 10'h090) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_215 = ((currYDiv == 10'h094) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_216 = ((currYDiv == 10'h098) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_217 = ((currYDiv == 10'h09c) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_218 = ((currYDiv == 10'h0a0) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_219 = ((currYDiv == 10'h0a4) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_220 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_221 = ((currYDiv == 10'h0ac) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_222 = ((currYDiv == 10'h0b0) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_223 = ((currYDiv == 10'h0b4) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_224 = ((currYDiv == 10'h0b8) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_225 = ((currYDiv == 10'h0bc) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_226 = ((currYDiv == 10'h0c0) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_227 = ((currYDiv == 10'h0c4) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_228 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_229 = ((currYDiv == 10'h0cc) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_230 = ((currYDiv == 10'h0d0) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_231 = ((currYDiv == 10'h0d4) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_232 = ((currYDiv == 10'h0d8) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_233 = ((currYDiv == 10'h0dc) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_234 = ((currYDiv == 10'h0e0) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_235 = ((currYDiv == 10'h0e4) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_236 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_237 = ((currYDiv == 10'h0ec) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_238 = ((currYDiv == 10'h0f0) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_239 = ((currYDiv == 10'h0f4) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_240 = ((currYDiv == 10'h0f8) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_241 = ((currYDiv == 10'h0fc) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_242 = ((currYDiv == 10'h100) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_243 = ((currYDiv == 10'h104) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_244 = ((currYDiv == 10'h108) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_245 = ((currYDiv == 10'h10c) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_246 = ((currYDiv == 10'h110) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_247 = ((currYDiv == 10'h114) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_248 = ((currYDiv == 10'h118) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_249 = ((currYDiv == 10'h11c) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_250 = ((currYDiv == 10'h120) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_251 = ((currYDiv == 10'h124) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l102_252 = ((currYDiv == 10'h02c) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_253 = ((currYDiv == 10'h030) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_254 = ((currYDiv == 10'h034) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_255 = ((currYDiv == 10'h038) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_256 = ((currYDiv == 10'h03c) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_257 = ((currYDiv == 10'h040) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_258 = ((currYDiv == 10'h044) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_259 = ((currYDiv == 10'h048) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_260 = ((currYDiv == 10'h04c) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_261 = ((currYDiv == 10'h050) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_262 = ((currYDiv == 10'h054) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_263 = ((currYDiv == 10'h058) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_264 = ((currYDiv == 10'h05c) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_265 = ((currYDiv == 10'h060) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_266 = ((currYDiv == 10'h064) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_267 = ((currYDiv == 10'h068) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_268 = ((currYDiv == 10'h06c) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_269 = ((currYDiv == 10'h070) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_270 = ((currYDiv == 10'h074) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_271 = ((currYDiv == 10'h078) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_272 = ((currYDiv == 10'h07c) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_273 = ((currYDiv == 10'h080) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_274 = ((currYDiv == 10'h084) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_275 = ((currYDiv == 10'h088) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_276 = ((currYDiv == 10'h08c) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_277 = ((currYDiv == 10'h090) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_278 = ((currYDiv == 10'h094) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_279 = ((currYDiv == 10'h098) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_280 = ((currYDiv == 10'h09c) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_281 = ((currYDiv == 10'h0a0) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_282 = ((currYDiv == 10'h0a4) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_283 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_284 = ((currYDiv == 10'h0ac) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_285 = ((currYDiv == 10'h0b0) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_286 = ((currYDiv == 10'h0b4) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_287 = ((currYDiv == 10'h0b8) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_288 = ((currYDiv == 10'h0bc) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_289 = ((currYDiv == 10'h0c0) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_290 = ((currYDiv == 10'h0c4) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_291 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_292 = ((currYDiv == 10'h0cc) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_293 = ((currYDiv == 10'h0d0) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_294 = ((currYDiv == 10'h0d4) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_295 = ((currYDiv == 10'h0d8) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_296 = ((currYDiv == 10'h0dc) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_297 = ((currYDiv == 10'h0e0) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_298 = ((currYDiv == 10'h0e4) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_299 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_300 = ((currYDiv == 10'h0ec) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_301 = ((currYDiv == 10'h0f0) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_302 = ((currYDiv == 10'h0f4) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_303 = ((currYDiv == 10'h0f8) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_304 = ((currYDiv == 10'h0fc) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_305 = ((currYDiv == 10'h100) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_306 = ((currYDiv == 10'h104) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_307 = ((currYDiv == 10'h108) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_308 = ((currYDiv == 10'h10c) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_309 = ((currYDiv == 10'h110) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_310 = ((currYDiv == 10'h114) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_311 = ((currYDiv == 10'h118) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_312 = ((currYDiv == 10'h11c) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_313 = ((currYDiv == 10'h120) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_314 = ((currYDiv == 10'h124) && (currXDiv == 10'h0fd));
  assign when_PictureGenerator_l102_315 = ((currYDiv == 10'h02c) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_316 = ((currYDiv == 10'h030) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_317 = ((currYDiv == 10'h034) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_318 = ((currYDiv == 10'h038) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_319 = ((currYDiv == 10'h03c) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_320 = ((currYDiv == 10'h040) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_321 = ((currYDiv == 10'h044) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_322 = ((currYDiv == 10'h048) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_323 = ((currYDiv == 10'h04c) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_324 = ((currYDiv == 10'h050) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_325 = ((currYDiv == 10'h054) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_326 = ((currYDiv == 10'h058) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_327 = ((currYDiv == 10'h05c) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_328 = ((currYDiv == 10'h060) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_329 = ((currYDiv == 10'h064) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_330 = ((currYDiv == 10'h068) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_331 = ((currYDiv == 10'h06c) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_332 = ((currYDiv == 10'h070) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_333 = ((currYDiv == 10'h074) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_334 = ((currYDiv == 10'h078) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_335 = ((currYDiv == 10'h07c) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_336 = ((currYDiv == 10'h080) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_337 = ((currYDiv == 10'h084) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_338 = ((currYDiv == 10'h088) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_339 = ((currYDiv == 10'h08c) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_340 = ((currYDiv == 10'h090) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_341 = ((currYDiv == 10'h094) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_342 = ((currYDiv == 10'h098) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_343 = ((currYDiv == 10'h09c) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_344 = ((currYDiv == 10'h0a0) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_345 = ((currYDiv == 10'h0a4) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_346 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_347 = ((currYDiv == 10'h0ac) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_348 = ((currYDiv == 10'h0b0) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_349 = ((currYDiv == 10'h0b4) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_350 = ((currYDiv == 10'h0b8) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_351 = ((currYDiv == 10'h0bc) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_352 = ((currYDiv == 10'h0c0) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_353 = ((currYDiv == 10'h0c4) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_354 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_355 = ((currYDiv == 10'h0cc) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_356 = ((currYDiv == 10'h0d0) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_357 = ((currYDiv == 10'h0d4) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_358 = ((currYDiv == 10'h0d8) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_359 = ((currYDiv == 10'h0dc) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_360 = ((currYDiv == 10'h0e0) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_361 = ((currYDiv == 10'h0e4) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_362 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_363 = ((currYDiv == 10'h0ec) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_364 = ((currYDiv == 10'h0f0) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_365 = ((currYDiv == 10'h0f4) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_366 = ((currYDiv == 10'h0f8) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_367 = ((currYDiv == 10'h0fc) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_368 = ((currYDiv == 10'h100) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_369 = ((currYDiv == 10'h104) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_370 = ((currYDiv == 10'h108) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_371 = ((currYDiv == 10'h10c) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_372 = ((currYDiv == 10'h110) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_373 = ((currYDiv == 10'h114) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_374 = ((currYDiv == 10'h118) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_375 = ((currYDiv == 10'h11c) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_376 = ((currYDiv == 10'h120) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_377 = ((currYDiv == 10'h124) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l102_378 = ((currYDiv == 10'h02c) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_379 = ((currYDiv == 10'h030) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_380 = ((currYDiv == 10'h034) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_381 = ((currYDiv == 10'h038) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_382 = ((currYDiv == 10'h03c) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_383 = ((currYDiv == 10'h040) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_384 = ((currYDiv == 10'h044) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_385 = ((currYDiv == 10'h048) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_386 = ((currYDiv == 10'h04c) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_387 = ((currYDiv == 10'h050) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_388 = ((currYDiv == 10'h054) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_389 = ((currYDiv == 10'h058) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_390 = ((currYDiv == 10'h05c) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_391 = ((currYDiv == 10'h060) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_392 = ((currYDiv == 10'h064) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_393 = ((currYDiv == 10'h068) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_394 = ((currYDiv == 10'h06c) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_395 = ((currYDiv == 10'h070) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_396 = ((currYDiv == 10'h074) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_397 = ((currYDiv == 10'h078) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_398 = ((currYDiv == 10'h07c) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_399 = ((currYDiv == 10'h080) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_400 = ((currYDiv == 10'h084) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_401 = ((currYDiv == 10'h088) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_402 = ((currYDiv == 10'h08c) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_403 = ((currYDiv == 10'h090) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_404 = ((currYDiv == 10'h094) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_405 = ((currYDiv == 10'h098) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_406 = ((currYDiv == 10'h09c) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_407 = ((currYDiv == 10'h0a0) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_408 = ((currYDiv == 10'h0a4) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_409 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_410 = ((currYDiv == 10'h0ac) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_411 = ((currYDiv == 10'h0b0) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_412 = ((currYDiv == 10'h0b4) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_413 = ((currYDiv == 10'h0b8) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_414 = ((currYDiv == 10'h0bc) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_415 = ((currYDiv == 10'h0c0) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_416 = ((currYDiv == 10'h0c4) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_417 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_418 = ((currYDiv == 10'h0cc) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_419 = ((currYDiv == 10'h0d0) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_420 = ((currYDiv == 10'h0d4) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_421 = ((currYDiv == 10'h0d8) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_422 = ((currYDiv == 10'h0dc) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_423 = ((currYDiv == 10'h0e0) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_424 = ((currYDiv == 10'h0e4) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_425 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_426 = ((currYDiv == 10'h0ec) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_427 = ((currYDiv == 10'h0f0) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_428 = ((currYDiv == 10'h0f4) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_429 = ((currYDiv == 10'h0f8) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_430 = ((currYDiv == 10'h0fc) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_431 = ((currYDiv == 10'h100) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_432 = ((currYDiv == 10'h104) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_433 = ((currYDiv == 10'h108) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_434 = ((currYDiv == 10'h10c) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_435 = ((currYDiv == 10'h110) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_436 = ((currYDiv == 10'h114) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_437 = ((currYDiv == 10'h118) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_438 = ((currYDiv == 10'h11c) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_439 = ((currYDiv == 10'h120) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_440 = ((currYDiv == 10'h124) && (currXDiv == 10'h139));
  assign when_PictureGenerator_l102_441 = ((currYDiv == 10'h02c) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_442 = ((currYDiv == 10'h030) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_443 = ((currYDiv == 10'h034) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_444 = ((currYDiv == 10'h038) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_445 = ((currYDiv == 10'h03c) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_446 = ((currYDiv == 10'h040) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_447 = ((currYDiv == 10'h044) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_448 = ((currYDiv == 10'h048) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_449 = ((currYDiv == 10'h04c) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_450 = ((currYDiv == 10'h050) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_451 = ((currYDiv == 10'h054) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_452 = ((currYDiv == 10'h058) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_453 = ((currYDiv == 10'h05c) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_454 = ((currYDiv == 10'h060) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_455 = ((currYDiv == 10'h064) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_456 = ((currYDiv == 10'h068) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_457 = ((currYDiv == 10'h06c) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_458 = ((currYDiv == 10'h070) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_459 = ((currYDiv == 10'h074) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_460 = ((currYDiv == 10'h078) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_461 = ((currYDiv == 10'h07c) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_462 = ((currYDiv == 10'h080) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_463 = ((currYDiv == 10'h084) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_464 = ((currYDiv == 10'h088) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_465 = ((currYDiv == 10'h08c) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_466 = ((currYDiv == 10'h090) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_467 = ((currYDiv == 10'h094) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_468 = ((currYDiv == 10'h098) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_469 = ((currYDiv == 10'h09c) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_470 = ((currYDiv == 10'h0a0) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_471 = ((currYDiv == 10'h0a4) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_472 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_473 = ((currYDiv == 10'h0ac) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_474 = ((currYDiv == 10'h0b0) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_475 = ((currYDiv == 10'h0b4) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_476 = ((currYDiv == 10'h0b8) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_477 = ((currYDiv == 10'h0bc) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_478 = ((currYDiv == 10'h0c0) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_479 = ((currYDiv == 10'h0c4) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_480 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_481 = ((currYDiv == 10'h0cc) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_482 = ((currYDiv == 10'h0d0) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_483 = ((currYDiv == 10'h0d4) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_484 = ((currYDiv == 10'h0d8) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_485 = ((currYDiv == 10'h0dc) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_486 = ((currYDiv == 10'h0e0) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_487 = ((currYDiv == 10'h0e4) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_488 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_489 = ((currYDiv == 10'h0ec) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_490 = ((currYDiv == 10'h0f0) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_491 = ((currYDiv == 10'h0f4) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_492 = ((currYDiv == 10'h0f8) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_493 = ((currYDiv == 10'h0fc) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_494 = ((currYDiv == 10'h100) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_495 = ((currYDiv == 10'h104) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_496 = ((currYDiv == 10'h108) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_497 = ((currYDiv == 10'h10c) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_498 = ((currYDiv == 10'h110) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_499 = ((currYDiv == 10'h114) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_500 = ((currYDiv == 10'h118) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_501 = ((currYDiv == 10'h11c) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_502 = ((currYDiv == 10'h120) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_503 = ((currYDiv == 10'h124) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l102_504 = ((currYDiv == 10'h02c) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_505 = ((currYDiv == 10'h030) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_506 = ((currYDiv == 10'h034) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_507 = ((currYDiv == 10'h038) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_508 = ((currYDiv == 10'h03c) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_509 = ((currYDiv == 10'h040) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_510 = ((currYDiv == 10'h044) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_511 = ((currYDiv == 10'h048) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_512 = ((currYDiv == 10'h04c) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_513 = ((currYDiv == 10'h050) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_514 = ((currYDiv == 10'h054) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_515 = ((currYDiv == 10'h058) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_516 = ((currYDiv == 10'h05c) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_517 = ((currYDiv == 10'h060) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_518 = ((currYDiv == 10'h064) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_519 = ((currYDiv == 10'h068) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_520 = ((currYDiv == 10'h06c) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_521 = ((currYDiv == 10'h070) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_522 = ((currYDiv == 10'h074) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_523 = ((currYDiv == 10'h078) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_524 = ((currYDiv == 10'h07c) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_525 = ((currYDiv == 10'h080) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_526 = ((currYDiv == 10'h084) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_527 = ((currYDiv == 10'h088) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_528 = ((currYDiv == 10'h08c) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_529 = ((currYDiv == 10'h090) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_530 = ((currYDiv == 10'h094) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_531 = ((currYDiv == 10'h098) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_532 = ((currYDiv == 10'h09c) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_533 = ((currYDiv == 10'h0a0) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_534 = ((currYDiv == 10'h0a4) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_535 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_536 = ((currYDiv == 10'h0ac) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_537 = ((currYDiv == 10'h0b0) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_538 = ((currYDiv == 10'h0b4) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_539 = ((currYDiv == 10'h0b8) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_540 = ((currYDiv == 10'h0bc) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_541 = ((currYDiv == 10'h0c0) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_542 = ((currYDiv == 10'h0c4) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_543 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_544 = ((currYDiv == 10'h0cc) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_545 = ((currYDiv == 10'h0d0) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_546 = ((currYDiv == 10'h0d4) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_547 = ((currYDiv == 10'h0d8) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_548 = ((currYDiv == 10'h0dc) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_549 = ((currYDiv == 10'h0e0) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_550 = ((currYDiv == 10'h0e4) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_551 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_552 = ((currYDiv == 10'h0ec) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_553 = ((currYDiv == 10'h0f0) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_554 = ((currYDiv == 10'h0f4) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_555 = ((currYDiv == 10'h0f8) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_556 = ((currYDiv == 10'h0fc) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_557 = ((currYDiv == 10'h100) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_558 = ((currYDiv == 10'h104) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_559 = ((currYDiv == 10'h108) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_560 = ((currYDiv == 10'h10c) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_561 = ((currYDiv == 10'h110) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_562 = ((currYDiv == 10'h114) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_563 = ((currYDiv == 10'h118) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_564 = ((currYDiv == 10'h11c) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_565 = ((currYDiv == 10'h120) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_566 = ((currYDiv == 10'h124) && (currXDiv == 10'h175));
  assign when_PictureGenerator_l102_567 = ((currYDiv == 10'h02c) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_568 = ((currYDiv == 10'h030) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_569 = ((currYDiv == 10'h034) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_570 = ((currYDiv == 10'h038) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_571 = ((currYDiv == 10'h03c) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_572 = ((currYDiv == 10'h040) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_573 = ((currYDiv == 10'h044) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_574 = ((currYDiv == 10'h048) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_575 = ((currYDiv == 10'h04c) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_576 = ((currYDiv == 10'h050) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_577 = ((currYDiv == 10'h054) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_578 = ((currYDiv == 10'h058) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_579 = ((currYDiv == 10'h05c) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_580 = ((currYDiv == 10'h060) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_581 = ((currYDiv == 10'h064) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_582 = ((currYDiv == 10'h068) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_583 = ((currYDiv == 10'h06c) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_584 = ((currYDiv == 10'h070) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_585 = ((currYDiv == 10'h074) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_586 = ((currYDiv == 10'h078) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_587 = ((currYDiv == 10'h07c) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_588 = ((currYDiv == 10'h080) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_589 = ((currYDiv == 10'h084) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_590 = ((currYDiv == 10'h088) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_591 = ((currYDiv == 10'h08c) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_592 = ((currYDiv == 10'h090) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_593 = ((currYDiv == 10'h094) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_594 = ((currYDiv == 10'h098) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_595 = ((currYDiv == 10'h09c) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_596 = ((currYDiv == 10'h0a0) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_597 = ((currYDiv == 10'h0a4) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_598 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_599 = ((currYDiv == 10'h0ac) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_600 = ((currYDiv == 10'h0b0) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_601 = ((currYDiv == 10'h0b4) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_602 = ((currYDiv == 10'h0b8) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_603 = ((currYDiv == 10'h0bc) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_604 = ((currYDiv == 10'h0c0) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_605 = ((currYDiv == 10'h0c4) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_606 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_607 = ((currYDiv == 10'h0cc) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_608 = ((currYDiv == 10'h0d0) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_609 = ((currYDiv == 10'h0d4) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_610 = ((currYDiv == 10'h0d8) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_611 = ((currYDiv == 10'h0dc) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_612 = ((currYDiv == 10'h0e0) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_613 = ((currYDiv == 10'h0e4) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_614 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_615 = ((currYDiv == 10'h0ec) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_616 = ((currYDiv == 10'h0f0) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_617 = ((currYDiv == 10'h0f4) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_618 = ((currYDiv == 10'h0f8) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_619 = ((currYDiv == 10'h0fc) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_620 = ((currYDiv == 10'h100) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_621 = ((currYDiv == 10'h104) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_622 = ((currYDiv == 10'h108) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_623 = ((currYDiv == 10'h10c) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_624 = ((currYDiv == 10'h110) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_625 = ((currYDiv == 10'h114) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_626 = ((currYDiv == 10'h118) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_627 = ((currYDiv == 10'h11c) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_628 = ((currYDiv == 10'h120) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l102_629 = ((currYDiv == 10'h124) && (currXDiv == 10'h193));
  assign when_PictureGenerator_l110 = ((currYDiv == 10'h048) && (currXDiv == 10'h06b));
  assign when_PictureGenerator_l110_1 = ((currYDiv == 10'h068) && (currXDiv == 10'h06b));
  assign when_PictureGenerator_l110_2 = ((currYDiv == 10'h088) && (currXDiv == 10'h06b));
  assign when_PictureGenerator_l110_3 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h06b));
  assign when_PictureGenerator_l110_4 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h06b));
  assign when_PictureGenerator_l110_5 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h06b));
  assign when_PictureGenerator_l110_6 = ((currYDiv == 10'h108) && (currXDiv == 10'h06b));
  assign when_PictureGenerator_l110_7 = ((currYDiv == 10'h048) && (currXDiv == 10'h06f));
  assign when_PictureGenerator_l110_8 = ((currYDiv == 10'h068) && (currXDiv == 10'h06f));
  assign when_PictureGenerator_l110_9 = ((currYDiv == 10'h088) && (currXDiv == 10'h06f));
  assign when_PictureGenerator_l110_10 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h06f));
  assign when_PictureGenerator_l110_11 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h06f));
  assign when_PictureGenerator_l110_12 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h06f));
  assign when_PictureGenerator_l110_13 = ((currYDiv == 10'h108) && (currXDiv == 10'h06f));
  assign when_PictureGenerator_l110_14 = ((currYDiv == 10'h048) && (currXDiv == 10'h073));
  assign when_PictureGenerator_l110_15 = ((currYDiv == 10'h068) && (currXDiv == 10'h073));
  assign when_PictureGenerator_l110_16 = ((currYDiv == 10'h088) && (currXDiv == 10'h073));
  assign when_PictureGenerator_l110_17 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h073));
  assign when_PictureGenerator_l110_18 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h073));
  assign when_PictureGenerator_l110_19 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h073));
  assign when_PictureGenerator_l110_20 = ((currYDiv == 10'h108) && (currXDiv == 10'h073));
  assign when_PictureGenerator_l110_21 = ((currYDiv == 10'h048) && (currXDiv == 10'h077));
  assign when_PictureGenerator_l110_22 = ((currYDiv == 10'h068) && (currXDiv == 10'h077));
  assign when_PictureGenerator_l110_23 = ((currYDiv == 10'h088) && (currXDiv == 10'h077));
  assign when_PictureGenerator_l110_24 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h077));
  assign when_PictureGenerator_l110_25 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h077));
  assign when_PictureGenerator_l110_26 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h077));
  assign when_PictureGenerator_l110_27 = ((currYDiv == 10'h108) && (currXDiv == 10'h077));
  assign when_PictureGenerator_l110_28 = ((currYDiv == 10'h048) && (currXDiv == 10'h07b));
  assign when_PictureGenerator_l110_29 = ((currYDiv == 10'h068) && (currXDiv == 10'h07b));
  assign when_PictureGenerator_l110_30 = ((currYDiv == 10'h088) && (currXDiv == 10'h07b));
  assign when_PictureGenerator_l110_31 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h07b));
  assign when_PictureGenerator_l110_32 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h07b));
  assign when_PictureGenerator_l110_33 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h07b));
  assign when_PictureGenerator_l110_34 = ((currYDiv == 10'h108) && (currXDiv == 10'h07b));
  assign when_PictureGenerator_l110_35 = ((currYDiv == 10'h048) && (currXDiv == 10'h07f));
  assign when_PictureGenerator_l110_36 = ((currYDiv == 10'h068) && (currXDiv == 10'h07f));
  assign when_PictureGenerator_l110_37 = ((currYDiv == 10'h088) && (currXDiv == 10'h07f));
  assign when_PictureGenerator_l110_38 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h07f));
  assign when_PictureGenerator_l110_39 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h07f));
  assign when_PictureGenerator_l110_40 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h07f));
  assign when_PictureGenerator_l110_41 = ((currYDiv == 10'h108) && (currXDiv == 10'h07f));
  assign when_PictureGenerator_l110_42 = ((currYDiv == 10'h048) && (currXDiv == 10'h083));
  assign when_PictureGenerator_l110_43 = ((currYDiv == 10'h068) && (currXDiv == 10'h083));
  assign when_PictureGenerator_l110_44 = ((currYDiv == 10'h088) && (currXDiv == 10'h083));
  assign when_PictureGenerator_l110_45 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h083));
  assign when_PictureGenerator_l110_46 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h083));
  assign when_PictureGenerator_l110_47 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h083));
  assign when_PictureGenerator_l110_48 = ((currYDiv == 10'h108) && (currXDiv == 10'h083));
  assign when_PictureGenerator_l110_49 = ((currYDiv == 10'h048) && (currXDiv == 10'h087));
  assign when_PictureGenerator_l110_50 = ((currYDiv == 10'h068) && (currXDiv == 10'h087));
  assign when_PictureGenerator_l110_51 = ((currYDiv == 10'h088) && (currXDiv == 10'h087));
  assign when_PictureGenerator_l110_52 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h087));
  assign when_PictureGenerator_l110_53 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h087));
  assign when_PictureGenerator_l110_54 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h087));
  assign when_PictureGenerator_l110_55 = ((currYDiv == 10'h108) && (currXDiv == 10'h087));
  assign when_PictureGenerator_l110_56 = ((currYDiv == 10'h048) && (currXDiv == 10'h08b));
  assign when_PictureGenerator_l110_57 = ((currYDiv == 10'h068) && (currXDiv == 10'h08b));
  assign when_PictureGenerator_l110_58 = ((currYDiv == 10'h088) && (currXDiv == 10'h08b));
  assign when_PictureGenerator_l110_59 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h08b));
  assign when_PictureGenerator_l110_60 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h08b));
  assign when_PictureGenerator_l110_61 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h08b));
  assign when_PictureGenerator_l110_62 = ((currYDiv == 10'h108) && (currXDiv == 10'h08b));
  assign when_PictureGenerator_l110_63 = ((currYDiv == 10'h048) && (currXDiv == 10'h08f));
  assign when_PictureGenerator_l110_64 = ((currYDiv == 10'h068) && (currXDiv == 10'h08f));
  assign when_PictureGenerator_l110_65 = ((currYDiv == 10'h088) && (currXDiv == 10'h08f));
  assign when_PictureGenerator_l110_66 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h08f));
  assign when_PictureGenerator_l110_67 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h08f));
  assign when_PictureGenerator_l110_68 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h08f));
  assign when_PictureGenerator_l110_69 = ((currYDiv == 10'h108) && (currXDiv == 10'h08f));
  assign when_PictureGenerator_l110_70 = ((currYDiv == 10'h048) && (currXDiv == 10'h093));
  assign when_PictureGenerator_l110_71 = ((currYDiv == 10'h068) && (currXDiv == 10'h093));
  assign when_PictureGenerator_l110_72 = ((currYDiv == 10'h088) && (currXDiv == 10'h093));
  assign when_PictureGenerator_l110_73 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h093));
  assign when_PictureGenerator_l110_74 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h093));
  assign when_PictureGenerator_l110_75 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h093));
  assign when_PictureGenerator_l110_76 = ((currYDiv == 10'h108) && (currXDiv == 10'h093));
  assign when_PictureGenerator_l110_77 = ((currYDiv == 10'h048) && (currXDiv == 10'h097));
  assign when_PictureGenerator_l110_78 = ((currYDiv == 10'h068) && (currXDiv == 10'h097));
  assign when_PictureGenerator_l110_79 = ((currYDiv == 10'h088) && (currXDiv == 10'h097));
  assign when_PictureGenerator_l110_80 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h097));
  assign when_PictureGenerator_l110_81 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h097));
  assign when_PictureGenerator_l110_82 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h097));
  assign when_PictureGenerator_l110_83 = ((currYDiv == 10'h108) && (currXDiv == 10'h097));
  assign when_PictureGenerator_l110_84 = ((currYDiv == 10'h048) && (currXDiv == 10'h09b));
  assign when_PictureGenerator_l110_85 = ((currYDiv == 10'h068) && (currXDiv == 10'h09b));
  assign when_PictureGenerator_l110_86 = ((currYDiv == 10'h088) && (currXDiv == 10'h09b));
  assign when_PictureGenerator_l110_87 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h09b));
  assign when_PictureGenerator_l110_88 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h09b));
  assign when_PictureGenerator_l110_89 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h09b));
  assign when_PictureGenerator_l110_90 = ((currYDiv == 10'h108) && (currXDiv == 10'h09b));
  assign when_PictureGenerator_l110_91 = ((currYDiv == 10'h048) && (currXDiv == 10'h09f));
  assign when_PictureGenerator_l110_92 = ((currYDiv == 10'h068) && (currXDiv == 10'h09f));
  assign when_PictureGenerator_l110_93 = ((currYDiv == 10'h088) && (currXDiv == 10'h09f));
  assign when_PictureGenerator_l110_94 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h09f));
  assign when_PictureGenerator_l110_95 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h09f));
  assign when_PictureGenerator_l110_96 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h09f));
  assign when_PictureGenerator_l110_97 = ((currYDiv == 10'h108) && (currXDiv == 10'h09f));
  assign when_PictureGenerator_l110_98 = ((currYDiv == 10'h048) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l110_99 = ((currYDiv == 10'h068) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l110_100 = ((currYDiv == 10'h088) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l110_101 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l110_102 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l110_103 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l110_104 = ((currYDiv == 10'h108) && (currXDiv == 10'h0a3));
  assign when_PictureGenerator_l110_105 = ((currYDiv == 10'h048) && (currXDiv == 10'h0a7));
  assign when_PictureGenerator_l110_106 = ((currYDiv == 10'h068) && (currXDiv == 10'h0a7));
  assign when_PictureGenerator_l110_107 = ((currYDiv == 10'h088) && (currXDiv == 10'h0a7));
  assign when_PictureGenerator_l110_108 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0a7));
  assign when_PictureGenerator_l110_109 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0a7));
  assign when_PictureGenerator_l110_110 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0a7));
  assign when_PictureGenerator_l110_111 = ((currYDiv == 10'h108) && (currXDiv == 10'h0a7));
  assign when_PictureGenerator_l110_112 = ((currYDiv == 10'h048) && (currXDiv == 10'h0ab));
  assign when_PictureGenerator_l110_113 = ((currYDiv == 10'h068) && (currXDiv == 10'h0ab));
  assign when_PictureGenerator_l110_114 = ((currYDiv == 10'h088) && (currXDiv == 10'h0ab));
  assign when_PictureGenerator_l110_115 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0ab));
  assign when_PictureGenerator_l110_116 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0ab));
  assign when_PictureGenerator_l110_117 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0ab));
  assign when_PictureGenerator_l110_118 = ((currYDiv == 10'h108) && (currXDiv == 10'h0ab));
  assign when_PictureGenerator_l110_119 = ((currYDiv == 10'h048) && (currXDiv == 10'h0af));
  assign when_PictureGenerator_l110_120 = ((currYDiv == 10'h068) && (currXDiv == 10'h0af));
  assign when_PictureGenerator_l110_121 = ((currYDiv == 10'h088) && (currXDiv == 10'h0af));
  assign when_PictureGenerator_l110_122 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0af));
  assign when_PictureGenerator_l110_123 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0af));
  assign when_PictureGenerator_l110_124 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0af));
  assign when_PictureGenerator_l110_125 = ((currYDiv == 10'h108) && (currXDiv == 10'h0af));
  assign when_PictureGenerator_l110_126 = ((currYDiv == 10'h048) && (currXDiv == 10'h0b3));
  assign when_PictureGenerator_l110_127 = ((currYDiv == 10'h068) && (currXDiv == 10'h0b3));
  assign when_PictureGenerator_l110_128 = ((currYDiv == 10'h088) && (currXDiv == 10'h0b3));
  assign when_PictureGenerator_l110_129 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0b3));
  assign when_PictureGenerator_l110_130 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0b3));
  assign when_PictureGenerator_l110_131 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0b3));
  assign when_PictureGenerator_l110_132 = ((currYDiv == 10'h108) && (currXDiv == 10'h0b3));
  assign when_PictureGenerator_l110_133 = ((currYDiv == 10'h048) && (currXDiv == 10'h0b7));
  assign when_PictureGenerator_l110_134 = ((currYDiv == 10'h068) && (currXDiv == 10'h0b7));
  assign when_PictureGenerator_l110_135 = ((currYDiv == 10'h088) && (currXDiv == 10'h0b7));
  assign when_PictureGenerator_l110_136 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0b7));
  assign when_PictureGenerator_l110_137 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0b7));
  assign when_PictureGenerator_l110_138 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0b7));
  assign when_PictureGenerator_l110_139 = ((currYDiv == 10'h108) && (currXDiv == 10'h0b7));
  assign when_PictureGenerator_l110_140 = ((currYDiv == 10'h048) && (currXDiv == 10'h0bb));
  assign when_PictureGenerator_l110_141 = ((currYDiv == 10'h068) && (currXDiv == 10'h0bb));
  assign when_PictureGenerator_l110_142 = ((currYDiv == 10'h088) && (currXDiv == 10'h0bb));
  assign when_PictureGenerator_l110_143 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0bb));
  assign when_PictureGenerator_l110_144 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0bb));
  assign when_PictureGenerator_l110_145 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0bb));
  assign when_PictureGenerator_l110_146 = ((currYDiv == 10'h108) && (currXDiv == 10'h0bb));
  assign when_PictureGenerator_l110_147 = ((currYDiv == 10'h048) && (currXDiv == 10'h0bf));
  assign when_PictureGenerator_l110_148 = ((currYDiv == 10'h068) && (currXDiv == 10'h0bf));
  assign when_PictureGenerator_l110_149 = ((currYDiv == 10'h088) && (currXDiv == 10'h0bf));
  assign when_PictureGenerator_l110_150 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0bf));
  assign when_PictureGenerator_l110_151 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0bf));
  assign when_PictureGenerator_l110_152 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0bf));
  assign when_PictureGenerator_l110_153 = ((currYDiv == 10'h108) && (currXDiv == 10'h0bf));
  assign when_PictureGenerator_l110_154 = ((currYDiv == 10'h048) && (currXDiv == 10'h0c3));
  assign when_PictureGenerator_l110_155 = ((currYDiv == 10'h068) && (currXDiv == 10'h0c3));
  assign when_PictureGenerator_l110_156 = ((currYDiv == 10'h088) && (currXDiv == 10'h0c3));
  assign when_PictureGenerator_l110_157 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0c3));
  assign when_PictureGenerator_l110_158 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0c3));
  assign when_PictureGenerator_l110_159 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0c3));
  assign when_PictureGenerator_l110_160 = ((currYDiv == 10'h108) && (currXDiv == 10'h0c3));
  assign when_PictureGenerator_l110_161 = ((currYDiv == 10'h048) && (currXDiv == 10'h0c7));
  assign when_PictureGenerator_l110_162 = ((currYDiv == 10'h068) && (currXDiv == 10'h0c7));
  assign when_PictureGenerator_l110_163 = ((currYDiv == 10'h088) && (currXDiv == 10'h0c7));
  assign when_PictureGenerator_l110_164 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0c7));
  assign when_PictureGenerator_l110_165 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0c7));
  assign when_PictureGenerator_l110_166 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0c7));
  assign when_PictureGenerator_l110_167 = ((currYDiv == 10'h108) && (currXDiv == 10'h0c7));
  assign when_PictureGenerator_l110_168 = ((currYDiv == 10'h048) && (currXDiv == 10'h0cb));
  assign when_PictureGenerator_l110_169 = ((currYDiv == 10'h068) && (currXDiv == 10'h0cb));
  assign when_PictureGenerator_l110_170 = ((currYDiv == 10'h088) && (currXDiv == 10'h0cb));
  assign when_PictureGenerator_l110_171 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0cb));
  assign when_PictureGenerator_l110_172 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0cb));
  assign when_PictureGenerator_l110_173 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0cb));
  assign when_PictureGenerator_l110_174 = ((currYDiv == 10'h108) && (currXDiv == 10'h0cb));
  assign when_PictureGenerator_l110_175 = ((currYDiv == 10'h048) && (currXDiv == 10'h0cf));
  assign when_PictureGenerator_l110_176 = ((currYDiv == 10'h068) && (currXDiv == 10'h0cf));
  assign when_PictureGenerator_l110_177 = ((currYDiv == 10'h088) && (currXDiv == 10'h0cf));
  assign when_PictureGenerator_l110_178 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0cf));
  assign when_PictureGenerator_l110_179 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0cf));
  assign when_PictureGenerator_l110_180 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0cf));
  assign when_PictureGenerator_l110_181 = ((currYDiv == 10'h108) && (currXDiv == 10'h0cf));
  assign when_PictureGenerator_l110_182 = ((currYDiv == 10'h048) && (currXDiv == 10'h0d3));
  assign when_PictureGenerator_l110_183 = ((currYDiv == 10'h068) && (currXDiv == 10'h0d3));
  assign when_PictureGenerator_l110_184 = ((currYDiv == 10'h088) && (currXDiv == 10'h0d3));
  assign when_PictureGenerator_l110_185 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0d3));
  assign when_PictureGenerator_l110_186 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0d3));
  assign when_PictureGenerator_l110_187 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0d3));
  assign when_PictureGenerator_l110_188 = ((currYDiv == 10'h108) && (currXDiv == 10'h0d3));
  assign when_PictureGenerator_l110_189 = ((currYDiv == 10'h048) && (currXDiv == 10'h0d7));
  assign when_PictureGenerator_l110_190 = ((currYDiv == 10'h068) && (currXDiv == 10'h0d7));
  assign when_PictureGenerator_l110_191 = ((currYDiv == 10'h088) && (currXDiv == 10'h0d7));
  assign when_PictureGenerator_l110_192 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0d7));
  assign when_PictureGenerator_l110_193 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0d7));
  assign when_PictureGenerator_l110_194 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0d7));
  assign when_PictureGenerator_l110_195 = ((currYDiv == 10'h108) && (currXDiv == 10'h0d7));
  assign when_PictureGenerator_l110_196 = ((currYDiv == 10'h048) && (currXDiv == 10'h0db));
  assign when_PictureGenerator_l110_197 = ((currYDiv == 10'h068) && (currXDiv == 10'h0db));
  assign when_PictureGenerator_l110_198 = ((currYDiv == 10'h088) && (currXDiv == 10'h0db));
  assign when_PictureGenerator_l110_199 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0db));
  assign when_PictureGenerator_l110_200 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0db));
  assign when_PictureGenerator_l110_201 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0db));
  assign when_PictureGenerator_l110_202 = ((currYDiv == 10'h108) && (currXDiv == 10'h0db));
  assign when_PictureGenerator_l110_203 = ((currYDiv == 10'h048) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l110_204 = ((currYDiv == 10'h068) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l110_205 = ((currYDiv == 10'h088) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l110_206 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l110_207 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l110_208 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l110_209 = ((currYDiv == 10'h108) && (currXDiv == 10'h0df));
  assign when_PictureGenerator_l110_210 = ((currYDiv == 10'h048) && (currXDiv == 10'h0e3));
  assign when_PictureGenerator_l110_211 = ((currYDiv == 10'h068) && (currXDiv == 10'h0e3));
  assign when_PictureGenerator_l110_212 = ((currYDiv == 10'h088) && (currXDiv == 10'h0e3));
  assign when_PictureGenerator_l110_213 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0e3));
  assign when_PictureGenerator_l110_214 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0e3));
  assign when_PictureGenerator_l110_215 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0e3));
  assign when_PictureGenerator_l110_216 = ((currYDiv == 10'h108) && (currXDiv == 10'h0e3));
  assign when_PictureGenerator_l110_217 = ((currYDiv == 10'h048) && (currXDiv == 10'h0e7));
  assign when_PictureGenerator_l110_218 = ((currYDiv == 10'h068) && (currXDiv == 10'h0e7));
  assign when_PictureGenerator_l110_219 = ((currYDiv == 10'h088) && (currXDiv == 10'h0e7));
  assign when_PictureGenerator_l110_220 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0e7));
  assign when_PictureGenerator_l110_221 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0e7));
  assign when_PictureGenerator_l110_222 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0e7));
  assign when_PictureGenerator_l110_223 = ((currYDiv == 10'h108) && (currXDiv == 10'h0e7));
  assign when_PictureGenerator_l110_224 = ((currYDiv == 10'h048) && (currXDiv == 10'h0eb));
  assign when_PictureGenerator_l110_225 = ((currYDiv == 10'h068) && (currXDiv == 10'h0eb));
  assign when_PictureGenerator_l110_226 = ((currYDiv == 10'h088) && (currXDiv == 10'h0eb));
  assign when_PictureGenerator_l110_227 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0eb));
  assign when_PictureGenerator_l110_228 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0eb));
  assign when_PictureGenerator_l110_229 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0eb));
  assign when_PictureGenerator_l110_230 = ((currYDiv == 10'h108) && (currXDiv == 10'h0eb));
  assign when_PictureGenerator_l110_231 = ((currYDiv == 10'h048) && (currXDiv == 10'h0ef));
  assign when_PictureGenerator_l110_232 = ((currYDiv == 10'h068) && (currXDiv == 10'h0ef));
  assign when_PictureGenerator_l110_233 = ((currYDiv == 10'h088) && (currXDiv == 10'h0ef));
  assign when_PictureGenerator_l110_234 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0ef));
  assign when_PictureGenerator_l110_235 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0ef));
  assign when_PictureGenerator_l110_236 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0ef));
  assign when_PictureGenerator_l110_237 = ((currYDiv == 10'h108) && (currXDiv == 10'h0ef));
  assign when_PictureGenerator_l110_238 = ((currYDiv == 10'h048) && (currXDiv == 10'h0f3));
  assign when_PictureGenerator_l110_239 = ((currYDiv == 10'h068) && (currXDiv == 10'h0f3));
  assign when_PictureGenerator_l110_240 = ((currYDiv == 10'h088) && (currXDiv == 10'h0f3));
  assign when_PictureGenerator_l110_241 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0f3));
  assign when_PictureGenerator_l110_242 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0f3));
  assign when_PictureGenerator_l110_243 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0f3));
  assign when_PictureGenerator_l110_244 = ((currYDiv == 10'h108) && (currXDiv == 10'h0f3));
  assign when_PictureGenerator_l110_245 = ((currYDiv == 10'h048) && (currXDiv == 10'h0f7));
  assign when_PictureGenerator_l110_246 = ((currYDiv == 10'h068) && (currXDiv == 10'h0f7));
  assign when_PictureGenerator_l110_247 = ((currYDiv == 10'h088) && (currXDiv == 10'h0f7));
  assign when_PictureGenerator_l110_248 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0f7));
  assign when_PictureGenerator_l110_249 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0f7));
  assign when_PictureGenerator_l110_250 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0f7));
  assign when_PictureGenerator_l110_251 = ((currYDiv == 10'h108) && (currXDiv == 10'h0f7));
  assign when_PictureGenerator_l110_252 = ((currYDiv == 10'h048) && (currXDiv == 10'h0fb));
  assign when_PictureGenerator_l110_253 = ((currYDiv == 10'h068) && (currXDiv == 10'h0fb));
  assign when_PictureGenerator_l110_254 = ((currYDiv == 10'h088) && (currXDiv == 10'h0fb));
  assign when_PictureGenerator_l110_255 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0fb));
  assign when_PictureGenerator_l110_256 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0fb));
  assign when_PictureGenerator_l110_257 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0fb));
  assign when_PictureGenerator_l110_258 = ((currYDiv == 10'h108) && (currXDiv == 10'h0fb));
  assign when_PictureGenerator_l110_259 = ((currYDiv == 10'h048) && (currXDiv == 10'h0ff));
  assign when_PictureGenerator_l110_260 = ((currYDiv == 10'h068) && (currXDiv == 10'h0ff));
  assign when_PictureGenerator_l110_261 = ((currYDiv == 10'h088) && (currXDiv == 10'h0ff));
  assign when_PictureGenerator_l110_262 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h0ff));
  assign when_PictureGenerator_l110_263 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h0ff));
  assign when_PictureGenerator_l110_264 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h0ff));
  assign when_PictureGenerator_l110_265 = ((currYDiv == 10'h108) && (currXDiv == 10'h0ff));
  assign when_PictureGenerator_l110_266 = ((currYDiv == 10'h048) && (currXDiv == 10'h103));
  assign when_PictureGenerator_l110_267 = ((currYDiv == 10'h068) && (currXDiv == 10'h103));
  assign when_PictureGenerator_l110_268 = ((currYDiv == 10'h088) && (currXDiv == 10'h103));
  assign when_PictureGenerator_l110_269 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h103));
  assign when_PictureGenerator_l110_270 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h103));
  assign when_PictureGenerator_l110_271 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h103));
  assign when_PictureGenerator_l110_272 = ((currYDiv == 10'h108) && (currXDiv == 10'h103));
  assign when_PictureGenerator_l110_273 = ((currYDiv == 10'h048) && (currXDiv == 10'h107));
  assign when_PictureGenerator_l110_274 = ((currYDiv == 10'h068) && (currXDiv == 10'h107));
  assign when_PictureGenerator_l110_275 = ((currYDiv == 10'h088) && (currXDiv == 10'h107));
  assign when_PictureGenerator_l110_276 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h107));
  assign when_PictureGenerator_l110_277 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h107));
  assign when_PictureGenerator_l110_278 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h107));
  assign when_PictureGenerator_l110_279 = ((currYDiv == 10'h108) && (currXDiv == 10'h107));
  assign when_PictureGenerator_l110_280 = ((currYDiv == 10'h048) && (currXDiv == 10'h10b));
  assign when_PictureGenerator_l110_281 = ((currYDiv == 10'h068) && (currXDiv == 10'h10b));
  assign when_PictureGenerator_l110_282 = ((currYDiv == 10'h088) && (currXDiv == 10'h10b));
  assign when_PictureGenerator_l110_283 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h10b));
  assign when_PictureGenerator_l110_284 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h10b));
  assign when_PictureGenerator_l110_285 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h10b));
  assign when_PictureGenerator_l110_286 = ((currYDiv == 10'h108) && (currXDiv == 10'h10b));
  assign when_PictureGenerator_l110_287 = ((currYDiv == 10'h048) && (currXDiv == 10'h10f));
  assign when_PictureGenerator_l110_288 = ((currYDiv == 10'h068) && (currXDiv == 10'h10f));
  assign when_PictureGenerator_l110_289 = ((currYDiv == 10'h088) && (currXDiv == 10'h10f));
  assign when_PictureGenerator_l110_290 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h10f));
  assign when_PictureGenerator_l110_291 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h10f));
  assign when_PictureGenerator_l110_292 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h10f));
  assign when_PictureGenerator_l110_293 = ((currYDiv == 10'h108) && (currXDiv == 10'h10f));
  assign when_PictureGenerator_l110_294 = ((currYDiv == 10'h048) && (currXDiv == 10'h113));
  assign when_PictureGenerator_l110_295 = ((currYDiv == 10'h068) && (currXDiv == 10'h113));
  assign when_PictureGenerator_l110_296 = ((currYDiv == 10'h088) && (currXDiv == 10'h113));
  assign when_PictureGenerator_l110_297 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h113));
  assign when_PictureGenerator_l110_298 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h113));
  assign when_PictureGenerator_l110_299 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h113));
  assign when_PictureGenerator_l110_300 = ((currYDiv == 10'h108) && (currXDiv == 10'h113));
  assign when_PictureGenerator_l110_301 = ((currYDiv == 10'h048) && (currXDiv == 10'h117));
  assign when_PictureGenerator_l110_302 = ((currYDiv == 10'h068) && (currXDiv == 10'h117));
  assign when_PictureGenerator_l110_303 = ((currYDiv == 10'h088) && (currXDiv == 10'h117));
  assign when_PictureGenerator_l110_304 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h117));
  assign when_PictureGenerator_l110_305 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h117));
  assign when_PictureGenerator_l110_306 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h117));
  assign when_PictureGenerator_l110_307 = ((currYDiv == 10'h108) && (currXDiv == 10'h117));
  assign when_PictureGenerator_l110_308 = ((currYDiv == 10'h048) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l110_309 = ((currYDiv == 10'h068) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l110_310 = ((currYDiv == 10'h088) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l110_311 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l110_312 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l110_313 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l110_314 = ((currYDiv == 10'h108) && (currXDiv == 10'h11b));
  assign when_PictureGenerator_l110_315 = ((currYDiv == 10'h048) && (currXDiv == 10'h11f));
  assign when_PictureGenerator_l110_316 = ((currYDiv == 10'h068) && (currXDiv == 10'h11f));
  assign when_PictureGenerator_l110_317 = ((currYDiv == 10'h088) && (currXDiv == 10'h11f));
  assign when_PictureGenerator_l110_318 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h11f));
  assign when_PictureGenerator_l110_319 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h11f));
  assign when_PictureGenerator_l110_320 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h11f));
  assign when_PictureGenerator_l110_321 = ((currYDiv == 10'h108) && (currXDiv == 10'h11f));
  assign when_PictureGenerator_l110_322 = ((currYDiv == 10'h048) && (currXDiv == 10'h123));
  assign when_PictureGenerator_l110_323 = ((currYDiv == 10'h068) && (currXDiv == 10'h123));
  assign when_PictureGenerator_l110_324 = ((currYDiv == 10'h088) && (currXDiv == 10'h123));
  assign when_PictureGenerator_l110_325 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h123));
  assign when_PictureGenerator_l110_326 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h123));
  assign when_PictureGenerator_l110_327 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h123));
  assign when_PictureGenerator_l110_328 = ((currYDiv == 10'h108) && (currXDiv == 10'h123));
  assign when_PictureGenerator_l110_329 = ((currYDiv == 10'h048) && (currXDiv == 10'h127));
  assign when_PictureGenerator_l110_330 = ((currYDiv == 10'h068) && (currXDiv == 10'h127));
  assign when_PictureGenerator_l110_331 = ((currYDiv == 10'h088) && (currXDiv == 10'h127));
  assign when_PictureGenerator_l110_332 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h127));
  assign when_PictureGenerator_l110_333 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h127));
  assign when_PictureGenerator_l110_334 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h127));
  assign when_PictureGenerator_l110_335 = ((currYDiv == 10'h108) && (currXDiv == 10'h127));
  assign when_PictureGenerator_l110_336 = ((currYDiv == 10'h048) && (currXDiv == 10'h12b));
  assign when_PictureGenerator_l110_337 = ((currYDiv == 10'h068) && (currXDiv == 10'h12b));
  assign when_PictureGenerator_l110_338 = ((currYDiv == 10'h088) && (currXDiv == 10'h12b));
  assign when_PictureGenerator_l110_339 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h12b));
  assign when_PictureGenerator_l110_340 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h12b));
  assign when_PictureGenerator_l110_341 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h12b));
  assign when_PictureGenerator_l110_342 = ((currYDiv == 10'h108) && (currXDiv == 10'h12b));
  assign when_PictureGenerator_l110_343 = ((currYDiv == 10'h048) && (currXDiv == 10'h12f));
  assign when_PictureGenerator_l110_344 = ((currYDiv == 10'h068) && (currXDiv == 10'h12f));
  assign when_PictureGenerator_l110_345 = ((currYDiv == 10'h088) && (currXDiv == 10'h12f));
  assign when_PictureGenerator_l110_346 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h12f));
  assign when_PictureGenerator_l110_347 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h12f));
  assign when_PictureGenerator_l110_348 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h12f));
  assign when_PictureGenerator_l110_349 = ((currYDiv == 10'h108) && (currXDiv == 10'h12f));
  assign when_PictureGenerator_l110_350 = ((currYDiv == 10'h048) && (currXDiv == 10'h133));
  assign when_PictureGenerator_l110_351 = ((currYDiv == 10'h068) && (currXDiv == 10'h133));
  assign when_PictureGenerator_l110_352 = ((currYDiv == 10'h088) && (currXDiv == 10'h133));
  assign when_PictureGenerator_l110_353 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h133));
  assign when_PictureGenerator_l110_354 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h133));
  assign when_PictureGenerator_l110_355 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h133));
  assign when_PictureGenerator_l110_356 = ((currYDiv == 10'h108) && (currXDiv == 10'h133));
  assign when_PictureGenerator_l110_357 = ((currYDiv == 10'h048) && (currXDiv == 10'h137));
  assign when_PictureGenerator_l110_358 = ((currYDiv == 10'h068) && (currXDiv == 10'h137));
  assign when_PictureGenerator_l110_359 = ((currYDiv == 10'h088) && (currXDiv == 10'h137));
  assign when_PictureGenerator_l110_360 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h137));
  assign when_PictureGenerator_l110_361 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h137));
  assign when_PictureGenerator_l110_362 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h137));
  assign when_PictureGenerator_l110_363 = ((currYDiv == 10'h108) && (currXDiv == 10'h137));
  assign when_PictureGenerator_l110_364 = ((currYDiv == 10'h048) && (currXDiv == 10'h13b));
  assign when_PictureGenerator_l110_365 = ((currYDiv == 10'h068) && (currXDiv == 10'h13b));
  assign when_PictureGenerator_l110_366 = ((currYDiv == 10'h088) && (currXDiv == 10'h13b));
  assign when_PictureGenerator_l110_367 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h13b));
  assign when_PictureGenerator_l110_368 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h13b));
  assign when_PictureGenerator_l110_369 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h13b));
  assign when_PictureGenerator_l110_370 = ((currYDiv == 10'h108) && (currXDiv == 10'h13b));
  assign when_PictureGenerator_l110_371 = ((currYDiv == 10'h048) && (currXDiv == 10'h13f));
  assign when_PictureGenerator_l110_372 = ((currYDiv == 10'h068) && (currXDiv == 10'h13f));
  assign when_PictureGenerator_l110_373 = ((currYDiv == 10'h088) && (currXDiv == 10'h13f));
  assign when_PictureGenerator_l110_374 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h13f));
  assign when_PictureGenerator_l110_375 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h13f));
  assign when_PictureGenerator_l110_376 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h13f));
  assign when_PictureGenerator_l110_377 = ((currYDiv == 10'h108) && (currXDiv == 10'h13f));
  assign when_PictureGenerator_l110_378 = ((currYDiv == 10'h048) && (currXDiv == 10'h143));
  assign when_PictureGenerator_l110_379 = ((currYDiv == 10'h068) && (currXDiv == 10'h143));
  assign when_PictureGenerator_l110_380 = ((currYDiv == 10'h088) && (currXDiv == 10'h143));
  assign when_PictureGenerator_l110_381 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h143));
  assign when_PictureGenerator_l110_382 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h143));
  assign when_PictureGenerator_l110_383 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h143));
  assign when_PictureGenerator_l110_384 = ((currYDiv == 10'h108) && (currXDiv == 10'h143));
  assign when_PictureGenerator_l110_385 = ((currYDiv == 10'h048) && (currXDiv == 10'h147));
  assign when_PictureGenerator_l110_386 = ((currYDiv == 10'h068) && (currXDiv == 10'h147));
  assign when_PictureGenerator_l110_387 = ((currYDiv == 10'h088) && (currXDiv == 10'h147));
  assign when_PictureGenerator_l110_388 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h147));
  assign when_PictureGenerator_l110_389 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h147));
  assign when_PictureGenerator_l110_390 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h147));
  assign when_PictureGenerator_l110_391 = ((currYDiv == 10'h108) && (currXDiv == 10'h147));
  assign when_PictureGenerator_l110_392 = ((currYDiv == 10'h048) && (currXDiv == 10'h14b));
  assign when_PictureGenerator_l110_393 = ((currYDiv == 10'h068) && (currXDiv == 10'h14b));
  assign when_PictureGenerator_l110_394 = ((currYDiv == 10'h088) && (currXDiv == 10'h14b));
  assign when_PictureGenerator_l110_395 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h14b));
  assign when_PictureGenerator_l110_396 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h14b));
  assign when_PictureGenerator_l110_397 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h14b));
  assign when_PictureGenerator_l110_398 = ((currYDiv == 10'h108) && (currXDiv == 10'h14b));
  assign when_PictureGenerator_l110_399 = ((currYDiv == 10'h048) && (currXDiv == 10'h14f));
  assign when_PictureGenerator_l110_400 = ((currYDiv == 10'h068) && (currXDiv == 10'h14f));
  assign when_PictureGenerator_l110_401 = ((currYDiv == 10'h088) && (currXDiv == 10'h14f));
  assign when_PictureGenerator_l110_402 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h14f));
  assign when_PictureGenerator_l110_403 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h14f));
  assign when_PictureGenerator_l110_404 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h14f));
  assign when_PictureGenerator_l110_405 = ((currYDiv == 10'h108) && (currXDiv == 10'h14f));
  assign when_PictureGenerator_l110_406 = ((currYDiv == 10'h048) && (currXDiv == 10'h153));
  assign when_PictureGenerator_l110_407 = ((currYDiv == 10'h068) && (currXDiv == 10'h153));
  assign when_PictureGenerator_l110_408 = ((currYDiv == 10'h088) && (currXDiv == 10'h153));
  assign when_PictureGenerator_l110_409 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h153));
  assign when_PictureGenerator_l110_410 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h153));
  assign when_PictureGenerator_l110_411 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h153));
  assign when_PictureGenerator_l110_412 = ((currYDiv == 10'h108) && (currXDiv == 10'h153));
  assign when_PictureGenerator_l110_413 = ((currYDiv == 10'h048) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l110_414 = ((currYDiv == 10'h068) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l110_415 = ((currYDiv == 10'h088) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l110_416 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l110_417 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l110_418 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l110_419 = ((currYDiv == 10'h108) && (currXDiv == 10'h157));
  assign when_PictureGenerator_l110_420 = ((currYDiv == 10'h048) && (currXDiv == 10'h15b));
  assign when_PictureGenerator_l110_421 = ((currYDiv == 10'h068) && (currXDiv == 10'h15b));
  assign when_PictureGenerator_l110_422 = ((currYDiv == 10'h088) && (currXDiv == 10'h15b));
  assign when_PictureGenerator_l110_423 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h15b));
  assign when_PictureGenerator_l110_424 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h15b));
  assign when_PictureGenerator_l110_425 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h15b));
  assign when_PictureGenerator_l110_426 = ((currYDiv == 10'h108) && (currXDiv == 10'h15b));
  assign when_PictureGenerator_l110_427 = ((currYDiv == 10'h048) && (currXDiv == 10'h15f));
  assign when_PictureGenerator_l110_428 = ((currYDiv == 10'h068) && (currXDiv == 10'h15f));
  assign when_PictureGenerator_l110_429 = ((currYDiv == 10'h088) && (currXDiv == 10'h15f));
  assign when_PictureGenerator_l110_430 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h15f));
  assign when_PictureGenerator_l110_431 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h15f));
  assign when_PictureGenerator_l110_432 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h15f));
  assign when_PictureGenerator_l110_433 = ((currYDiv == 10'h108) && (currXDiv == 10'h15f));
  assign when_PictureGenerator_l110_434 = ((currYDiv == 10'h048) && (currXDiv == 10'h163));
  assign when_PictureGenerator_l110_435 = ((currYDiv == 10'h068) && (currXDiv == 10'h163));
  assign when_PictureGenerator_l110_436 = ((currYDiv == 10'h088) && (currXDiv == 10'h163));
  assign when_PictureGenerator_l110_437 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h163));
  assign when_PictureGenerator_l110_438 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h163));
  assign when_PictureGenerator_l110_439 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h163));
  assign when_PictureGenerator_l110_440 = ((currYDiv == 10'h108) && (currXDiv == 10'h163));
  assign when_PictureGenerator_l110_441 = ((currYDiv == 10'h048) && (currXDiv == 10'h167));
  assign when_PictureGenerator_l110_442 = ((currYDiv == 10'h068) && (currXDiv == 10'h167));
  assign when_PictureGenerator_l110_443 = ((currYDiv == 10'h088) && (currXDiv == 10'h167));
  assign when_PictureGenerator_l110_444 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h167));
  assign when_PictureGenerator_l110_445 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h167));
  assign when_PictureGenerator_l110_446 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h167));
  assign when_PictureGenerator_l110_447 = ((currYDiv == 10'h108) && (currXDiv == 10'h167));
  assign when_PictureGenerator_l110_448 = ((currYDiv == 10'h048) && (currXDiv == 10'h16b));
  assign when_PictureGenerator_l110_449 = ((currYDiv == 10'h068) && (currXDiv == 10'h16b));
  assign when_PictureGenerator_l110_450 = ((currYDiv == 10'h088) && (currXDiv == 10'h16b));
  assign when_PictureGenerator_l110_451 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h16b));
  assign when_PictureGenerator_l110_452 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h16b));
  assign when_PictureGenerator_l110_453 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h16b));
  assign when_PictureGenerator_l110_454 = ((currYDiv == 10'h108) && (currXDiv == 10'h16b));
  assign when_PictureGenerator_l110_455 = ((currYDiv == 10'h048) && (currXDiv == 10'h16f));
  assign when_PictureGenerator_l110_456 = ((currYDiv == 10'h068) && (currXDiv == 10'h16f));
  assign when_PictureGenerator_l110_457 = ((currYDiv == 10'h088) && (currXDiv == 10'h16f));
  assign when_PictureGenerator_l110_458 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h16f));
  assign when_PictureGenerator_l110_459 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h16f));
  assign when_PictureGenerator_l110_460 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h16f));
  assign when_PictureGenerator_l110_461 = ((currYDiv == 10'h108) && (currXDiv == 10'h16f));
  assign when_PictureGenerator_l110_462 = ((currYDiv == 10'h048) && (currXDiv == 10'h173));
  assign when_PictureGenerator_l110_463 = ((currYDiv == 10'h068) && (currXDiv == 10'h173));
  assign when_PictureGenerator_l110_464 = ((currYDiv == 10'h088) && (currXDiv == 10'h173));
  assign when_PictureGenerator_l110_465 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h173));
  assign when_PictureGenerator_l110_466 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h173));
  assign when_PictureGenerator_l110_467 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h173));
  assign when_PictureGenerator_l110_468 = ((currYDiv == 10'h108) && (currXDiv == 10'h173));
  assign when_PictureGenerator_l110_469 = ((currYDiv == 10'h048) && (currXDiv == 10'h177));
  assign when_PictureGenerator_l110_470 = ((currYDiv == 10'h068) && (currXDiv == 10'h177));
  assign when_PictureGenerator_l110_471 = ((currYDiv == 10'h088) && (currXDiv == 10'h177));
  assign when_PictureGenerator_l110_472 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h177));
  assign when_PictureGenerator_l110_473 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h177));
  assign when_PictureGenerator_l110_474 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h177));
  assign when_PictureGenerator_l110_475 = ((currYDiv == 10'h108) && (currXDiv == 10'h177));
  assign when_PictureGenerator_l110_476 = ((currYDiv == 10'h048) && (currXDiv == 10'h17b));
  assign when_PictureGenerator_l110_477 = ((currYDiv == 10'h068) && (currXDiv == 10'h17b));
  assign when_PictureGenerator_l110_478 = ((currYDiv == 10'h088) && (currXDiv == 10'h17b));
  assign when_PictureGenerator_l110_479 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h17b));
  assign when_PictureGenerator_l110_480 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h17b));
  assign when_PictureGenerator_l110_481 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h17b));
  assign when_PictureGenerator_l110_482 = ((currYDiv == 10'h108) && (currXDiv == 10'h17b));
  assign when_PictureGenerator_l110_483 = ((currYDiv == 10'h048) && (currXDiv == 10'h17f));
  assign when_PictureGenerator_l110_484 = ((currYDiv == 10'h068) && (currXDiv == 10'h17f));
  assign when_PictureGenerator_l110_485 = ((currYDiv == 10'h088) && (currXDiv == 10'h17f));
  assign when_PictureGenerator_l110_486 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h17f));
  assign when_PictureGenerator_l110_487 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h17f));
  assign when_PictureGenerator_l110_488 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h17f));
  assign when_PictureGenerator_l110_489 = ((currYDiv == 10'h108) && (currXDiv == 10'h17f));
  assign when_PictureGenerator_l110_490 = ((currYDiv == 10'h048) && (currXDiv == 10'h183));
  assign when_PictureGenerator_l110_491 = ((currYDiv == 10'h068) && (currXDiv == 10'h183));
  assign when_PictureGenerator_l110_492 = ((currYDiv == 10'h088) && (currXDiv == 10'h183));
  assign when_PictureGenerator_l110_493 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h183));
  assign when_PictureGenerator_l110_494 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h183));
  assign when_PictureGenerator_l110_495 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h183));
  assign when_PictureGenerator_l110_496 = ((currYDiv == 10'h108) && (currXDiv == 10'h183));
  assign when_PictureGenerator_l110_497 = ((currYDiv == 10'h048) && (currXDiv == 10'h187));
  assign when_PictureGenerator_l110_498 = ((currYDiv == 10'h068) && (currXDiv == 10'h187));
  assign when_PictureGenerator_l110_499 = ((currYDiv == 10'h088) && (currXDiv == 10'h187));
  assign when_PictureGenerator_l110_500 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h187));
  assign when_PictureGenerator_l110_501 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h187));
  assign when_PictureGenerator_l110_502 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h187));
  assign when_PictureGenerator_l110_503 = ((currYDiv == 10'h108) && (currXDiv == 10'h187));
  assign when_PictureGenerator_l110_504 = ((currYDiv == 10'h048) && (currXDiv == 10'h18b));
  assign when_PictureGenerator_l110_505 = ((currYDiv == 10'h068) && (currXDiv == 10'h18b));
  assign when_PictureGenerator_l110_506 = ((currYDiv == 10'h088) && (currXDiv == 10'h18b));
  assign when_PictureGenerator_l110_507 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h18b));
  assign when_PictureGenerator_l110_508 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h18b));
  assign when_PictureGenerator_l110_509 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h18b));
  assign when_PictureGenerator_l110_510 = ((currYDiv == 10'h108) && (currXDiv == 10'h18b));
  assign when_PictureGenerator_l110_511 = ((currYDiv == 10'h048) && (currXDiv == 10'h18f));
  assign when_PictureGenerator_l110_512 = ((currYDiv == 10'h068) && (currXDiv == 10'h18f));
  assign when_PictureGenerator_l110_513 = ((currYDiv == 10'h088) && (currXDiv == 10'h18f));
  assign when_PictureGenerator_l110_514 = ((currYDiv == 10'h0a8) && (currXDiv == 10'h18f));
  assign when_PictureGenerator_l110_515 = ((currYDiv == 10'h0c8) && (currXDiv == 10'h18f));
  assign when_PictureGenerator_l110_516 = ((currYDiv == 10'h0e8) && (currXDiv == 10'h18f));
  assign when_PictureGenerator_l110_517 = ((currYDiv == 10'h108) && (currXDiv == 10'h18f));
  assign when_PictureGenerator_l115 = ((((currYDiv == 10'h027) || (currYDiv == 10'h129)) && (10'h069 <= currXDiv)) && (currXDiv <= 10'h193));
  assign when_PictureGenerator_l117 = (((10'h027 <= currYDiv) && (currYDiv <= 10'h129)) && ((currXDiv == 10'h069) || (currXDiv == 10'h193)));
  assign when_PictureGenerator_l119 = (((((10'h067 < currXDiv) && (currXDiv < 10'h193)) && (10'h027 < currYDiv)) && (currYDiv < 10'h128)) && (16'h0000 < colorInRam));
  assign when_PictureGenerator_l121 = (((currYDiv == 10'h0a8) && (10'h068 < currXDiv)) && (currXDiv <= 10'h193));
  assign ram_addr = rAddr_ram_addr;
  always @(*) begin
    rAddr_ram_x = 10'h000;
    if(when_PictureGenerator_l130) begin
      rAddr_ram_x = (currXDiv - 10'h068);
    end
  end

  always @(*) begin
    rAddr_ram_y = 10'h000;
    if(when_PictureGenerator_l130) begin
      rAddr_ram_y = (currYDiv - 10'h028);
    end
  end

  always @(*) begin
    ram_en = rAddr_ram_en;
    if(!when_PictureGenerator_l130) begin
      ram_en = 5'h00;
    end
  end

  assign when_PictureGenerator_l130 = ((((10'h067 < currXDiv) && (currXDiv < 10'h194)) && (10'h027 < currYDiv)) && (currYDiv < 10'h128));
  assign _zz_when_PictureGenerator_l78 = 12'h19a;
  assign _zz_when_PictureGenerator_l87 = 12'h00f;
  always @(*) begin
    _zz_when_PictureGenerator_l138_1 = _zz__zz_when_PictureGenerator_l138_1[7:0];
    if(when_PictureGenerator_l78) begin
      _zz_when_PictureGenerator_l138_1 = _zz__zz_when_PictureGenerator_l138_1_3[7:0];
    end else begin
      if(when_PictureGenerator_l81) begin
        _zz_when_PictureGenerator_l138_1 = _zz__zz_when_PictureGenerator_l138_1_6[7:0];
      end
    end
  end

  always @(*) begin
    _zz_when_PictureGenerator_l138 = _zz__zz_when_PictureGenerator_l138;
    if(when_PictureGenerator_l78) begin
      _zz_when_PictureGenerator_l138 = _zz__zz_when_PictureGenerator_l138_9;
    end else begin
      if(when_PictureGenerator_l81) begin
        _zz_when_PictureGenerator_l138 = _zz__zz_when_PictureGenerator_l138_18;
      end
    end
  end

  assign when_PictureGenerator_l78 = (_zz_when_PictureGenerator_l78_5 < _zz_when_PictureGenerator_l78_6);
  assign when_PictureGenerator_l81 = (_zz_when_PictureGenerator_l81 < _zz_when_PictureGenerator_l81_1);
  assign when_PictureGenerator_l87 = ((((_zz_when_PictureGenerator_l78 <= _zz_when_PictureGenerator_l87_5) && (_zz_when_PictureGenerator_l87 <= _zz_when_PictureGenerator_l87_6)) && (_zz_when_PictureGenerator_l87_7 < _zz_when_PictureGenerator_l87_8)) && (_zz_when_PictureGenerator_l87_9 < _zz_when_PictureGenerator_l87_10));
  always @(*) begin
    if(when_PictureGenerator_l87) begin
      when_PictureGenerator_l138 = _zz_when_PictureGenerator_l138[_zz_when_PictureGenerator_l138_10];
    end else begin
      when_PictureGenerator_l138 = 1'b0;
    end
  end

  assign _zz_when_PictureGenerator_l78_1 = 12'h1b2;
  assign _zz_when_PictureGenerator_l87_1 = 12'h00f;
  always @(*) begin
    _zz_when_PictureGenerator_l138_3 = _zz__zz_when_PictureGenerator_l138_3_1[7:0];
    if(when_PictureGenerator_l78_1) begin
      _zz_when_PictureGenerator_l138_3 = _zz__zz_when_PictureGenerator_l138_3_4[7:0];
    end else begin
      if(when_PictureGenerator_l81_1) begin
        _zz_when_PictureGenerator_l138_3 = _zz__zz_when_PictureGenerator_l138_3_7[7:0];
      end
    end
  end

  always @(*) begin
    _zz_when_PictureGenerator_l138_2 = _zz__zz_when_PictureGenerator_l138_2_1;
    if(when_PictureGenerator_l78_1) begin
      _zz_when_PictureGenerator_l138_2 = _zz__zz_when_PictureGenerator_l138_2_9;
    end else begin
      if(when_PictureGenerator_l81_1) begin
        _zz_when_PictureGenerator_l138_2 = _zz__zz_when_PictureGenerator_l138_2_18;
      end
    end
  end

  assign when_PictureGenerator_l78_1 = (_zz_when_PictureGenerator_l78_1_1 < _zz_when_PictureGenerator_l78_1_2);
  assign when_PictureGenerator_l81_1 = (_zz_when_PictureGenerator_l81_1_1 < _zz_when_PictureGenerator_l81_1_2);
  assign when_PictureGenerator_l87_1 = ((((_zz_when_PictureGenerator_l78_1 <= _zz_when_PictureGenerator_l87_1_1) && (_zz_when_PictureGenerator_l87_1 <= _zz_when_PictureGenerator_l87_1_2)) && (_zz_when_PictureGenerator_l87_1_3 < _zz_when_PictureGenerator_l87_1_4)) && (_zz_when_PictureGenerator_l87_1_5 < _zz_when_PictureGenerator_l87_1_6));
  always @(*) begin
    if(when_PictureGenerator_l87_1) begin
      when_PictureGenerator_l138_1 = _zz_when_PictureGenerator_l138_2[_zz_when_PictureGenerator_l138_1_1];
    end else begin
      when_PictureGenerator_l138_1 = 1'b0;
    end
  end

  assign _zz_when_PictureGenerator_l78_2 = 12'h1ca;
  assign _zz_when_PictureGenerator_l87_2 = 12'h00f;
  always @(*) begin
    _zz_when_PictureGenerator_l138_5 = _zz__zz_when_PictureGenerator_l138_5_1[7:0];
    if(when_PictureGenerator_l78_2) begin
      _zz_when_PictureGenerator_l138_5 = _zz__zz_when_PictureGenerator_l138_5_4[7:0];
    end else begin
      if(when_PictureGenerator_l81_2) begin
        _zz_when_PictureGenerator_l138_5 = _zz__zz_when_PictureGenerator_l138_5_7[7:0];
      end
    end
  end

  always @(*) begin
    _zz_when_PictureGenerator_l138_4 = _zz__zz_when_PictureGenerator_l138_4_1;
    if(when_PictureGenerator_l78_2) begin
      _zz_when_PictureGenerator_l138_4 = _zz__zz_when_PictureGenerator_l138_4_9;
    end else begin
      if(when_PictureGenerator_l81_2) begin
        _zz_when_PictureGenerator_l138_4 = _zz__zz_when_PictureGenerator_l138_4_18;
      end
    end
  end

  assign when_PictureGenerator_l78_2 = (_zz_when_PictureGenerator_l78_2_1 < _zz_when_PictureGenerator_l78_2_2);
  assign when_PictureGenerator_l81_2 = (_zz_when_PictureGenerator_l81_2 < _zz_when_PictureGenerator_l81_2_1);
  assign when_PictureGenerator_l87_2 = ((((_zz_when_PictureGenerator_l78_2 <= _zz_when_PictureGenerator_l87_2_1) && (_zz_when_PictureGenerator_l87_2 <= _zz_when_PictureGenerator_l87_2_2)) && (_zz_when_PictureGenerator_l87_2_3 < _zz_when_PictureGenerator_l87_2_4)) && (_zz_when_PictureGenerator_l87_2_5 < _zz_when_PictureGenerator_l87_2_6));
  always @(*) begin
    if(when_PictureGenerator_l87_2) begin
      when_PictureGenerator_l138_2 = _zz_when_PictureGenerator_l138_4[_zz_when_PictureGenerator_l138_2_1];
    end else begin
      when_PictureGenerator_l138_2 = 1'b0;
    end
  end

  assign _zz_when_PictureGenerator_l78_3 = 12'h1e2;
  assign _zz_when_PictureGenerator_l87_3 = 12'h00f;
  always @(*) begin
    _zz_when_PictureGenerator_l138_7 = _zz__zz_when_PictureGenerator_l138_7_1[7:0];
    if(when_PictureGenerator_l78_3) begin
      _zz_when_PictureGenerator_l138_7 = _zz__zz_when_PictureGenerator_l138_7_4[7:0];
    end else begin
      if(when_PictureGenerator_l81_3) begin
        _zz_when_PictureGenerator_l138_7 = _zz__zz_when_PictureGenerator_l138_7_7[7:0];
      end
    end
  end

  always @(*) begin
    _zz_when_PictureGenerator_l138_6 = _zz__zz_when_PictureGenerator_l138_6_1;
    if(when_PictureGenerator_l78_3) begin
      _zz_when_PictureGenerator_l138_6 = _zz__zz_when_PictureGenerator_l138_6_9;
    end else begin
      if(when_PictureGenerator_l81_3) begin
        _zz_when_PictureGenerator_l138_6 = _zz__zz_when_PictureGenerator_l138_6_18;
      end
    end
  end

  assign when_PictureGenerator_l78_3 = (_zz_when_PictureGenerator_l78_3_1 < _zz_when_PictureGenerator_l78_3_2);
  assign when_PictureGenerator_l81_3 = (_zz_when_PictureGenerator_l81_3 < _zz_when_PictureGenerator_l81_3_1);
  assign when_PictureGenerator_l87_3 = ((((_zz_when_PictureGenerator_l78_3 <= _zz_when_PictureGenerator_l87_3_1) && (_zz_when_PictureGenerator_l87_3 <= _zz_when_PictureGenerator_l87_3_2)) && (_zz_when_PictureGenerator_l87_3_3 < _zz_when_PictureGenerator_l87_3_4)) && (_zz_when_PictureGenerator_l87_3_5 < _zz_when_PictureGenerator_l87_3_6));
  always @(*) begin
    if(when_PictureGenerator_l87_3) begin
      when_PictureGenerator_l138_3 = _zz_when_PictureGenerator_l138_6[_zz_when_PictureGenerator_l138_3_1];
    end else begin
      when_PictureGenerator_l138_3 = 1'b0;
    end
  end

  assign _zz_when_PictureGenerator_l78_4 = 12'h1fa;
  assign _zz_when_PictureGenerator_l87_4 = 12'h00f;
  always @(*) begin
    _zz_when_PictureGenerator_l138_9 = _zz__zz_when_PictureGenerator_l138_9_1[7:0];
    if(when_PictureGenerator_l78_4) begin
      _zz_when_PictureGenerator_l138_9 = _zz__zz_when_PictureGenerator_l138_9_4[7:0];
    end else begin
      if(when_PictureGenerator_l81_4) begin
        _zz_when_PictureGenerator_l138_9 = _zz__zz_when_PictureGenerator_l138_9_7[7:0];
      end
    end
  end

  always @(*) begin
    _zz_when_PictureGenerator_l138_8 = _zz__zz_when_PictureGenerator_l138_8_1;
    if(when_PictureGenerator_l78_4) begin
      _zz_when_PictureGenerator_l138_8 = _zz__zz_when_PictureGenerator_l138_8_9;
    end else begin
      if(when_PictureGenerator_l81_4) begin
        _zz_when_PictureGenerator_l138_8 = _zz__zz_when_PictureGenerator_l138_8_18;
      end
    end
  end

  assign when_PictureGenerator_l78_4 = (_zz_when_PictureGenerator_l78_4_1 < _zz_when_PictureGenerator_l78_4_2);
  assign when_PictureGenerator_l81_4 = (_zz_when_PictureGenerator_l81_4 < _zz_when_PictureGenerator_l81_4_1);
  assign when_PictureGenerator_l87_4 = ((((_zz_when_PictureGenerator_l78_4 <= _zz_when_PictureGenerator_l87_4_1) && (_zz_when_PictureGenerator_l87_4 <= _zz_when_PictureGenerator_l87_4_2)) && (_zz_when_PictureGenerator_l87_4_3 < _zz_when_PictureGenerator_l87_4_4)) && (_zz_when_PictureGenerator_l87_4_5 < _zz_when_PictureGenerator_l87_4_6));
  always @(*) begin
    if(when_PictureGenerator_l87_4) begin
      when_PictureGenerator_l138_4 = _zz_when_PictureGenerator_l138_8[_zz_when_PictureGenerator_l138_4_1];
    end else begin
      when_PictureGenerator_l138_4 = 1'b0;
    end
  end

  always @(posedge clk or posedge reset) begin
    if(reset) begin
      colorInRam <= 16'h0000;
    end else begin
      colorInRam <= ram_color;
    end
  end


endmodule

module RAddressGen (
  output     [4:0]    ram_en,
  input      [9:0]    ram_x,
  input      [9:0]    ram_y,
  output     [13:0]   ram_addr,
  input               clk,
  input               reset
);

  wire       [7:0]    _zz_ram_addr;
  wire       [5:0]    _zz_ram_addr_1;
  wire       [13:0]   _zz_ram_addr_2;
  wire       [0:0]    _zz_ram_addr_3;
  wire       [2:0]    filmSel;
  reg        [4:0]    en;
  wire       [2:0]    switch_AddressGen_l27;

  assign _zz_ram_addr = ram_y[7:0];
  assign _zz_ram_addr_1 = ram_x[5:0];
  assign _zz_ram_addr_3 = 1'b0;
  assign _zz_ram_addr_2 = {13'd0, _zz_ram_addr_3};
  assign filmSel = {{ram_x[8],ram_x[7]},ram_x[6]};
  assign switch_AddressGen_l27 = filmSel;
  assign ram_en = en;
  assign ram_addr = ((|ram_en) ? {_zz_ram_addr,_zz_ram_addr_1} : _zz_ram_addr_2);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      en <= 5'h00;
    end else begin
      case(switch_AddressGen_l27)
        3'b000 : begin
          en <= 5'h01;
        end
        3'b001 : begin
          en <= 5'h02;
        end
        3'b010 : begin
          en <= 5'h04;
        end
        3'b011 : begin
          en <= 5'h08;
        end
        default : begin
          en <= 5'h10;
        end
      endcase
    end
  end


endmodule
